PK   G��X� �pO#  	B    cirkitFile.json���ȕ�o�P`h:u��/3I�vf�L��aE�ڴ��Z=�Y��7�״uȶ[-J�b��l��vc[b�zxT:U/�:�q�m~���lc�S�ެ6��%��Żf�}h�_5��պ�m�������G�w���:f�ml��&��mh��4}�Ă2�*[Ʀɺ�i�i\��mmj��|����
$V05��
��b�����A�`j/f�*�:��
���RSb���K1�T�ԕ�A��r�<Q�% U�s%ɓ�X"Q�ӥX"Q��X"Q�S�X"Qȓ�X"Q��� q/�n�_o�q��������Yӆ>�eo�j�����]YtE�sk�ȓ� ��3����){�x�x�	Xy�$���ȇ�A��?i'��9���A���|�K$
�%�H�J,�(�#�X"Q�G(�D���2b	�C��B>�w�t�d�^:gp�t/�H�-�H�)���yW,�(�yW,�(�yW,�(�yW,�(�yW,�(�yW,aj/ϻb�D!ϝb�D!ϝb�D!ϝb�D�-ϝ^�;��B�;��B�;��B�;��B�;����)�H��)�H��)�H��)�H��)�H��x���S,�(�S,�(�S,�(�S,a�\�;��B�;��B�;'כq�m����ϡ�כ�f����� ���G�a�Kg� 4v�����t����Yl�t��3����ac�#,]���yl�t��Ksl�6vP:�ҥ��;(a�L]`cW`c�#,��Kl�Jl�t��3u��]�����t��&xrvX>��������^�������|��/8~`���#0?���i`���OV��vX>��3�������|�4;8~`ׁ�#0?K��y`���O��vX>��B�f�������1���X>��"
p��w8з8��Â���,��x�	8~`���#0����?�|��?�������|�V	?������WY���X>���0p����G`>^�~H�?�|��uu�������|�"?�������2��~�
���8��p`���#0���?�|�㕯�������|�f?������W���X>��:ip����G`>^ፍ��,��xm:8~`���#0����?�|��z �������|\� ?�J�R���`�����G`>���`���u/���,���b8~`���#0���?�|��*)��������뻀��X>�qep����G`>����`���Հ���,����8~������`���#�����|\;
?�������^���X>�q�.p����G`>�4��_�X>�q�4p����G`>����`��	��U�K���E������懕Dg������|z~���O?,�9��a�Ι��l�l~Xsn��vza���7����Ovc����j�����w�wٳ6?�|���l���M�$9�H?ވ>^:d<����x&[<�m/��X��ɾ~��J<��+�q���D��+[4���!��w���K>k}��.�J��G�kg5~���Y�O��:WUmX6Y��ͼ5MV���F�e�ۼ����Y�O�{H�:��b:oh��>��E��,����M��j.��ӑ�E�U��YYR�y�����vI�]V�R��Y���bWfI&d��L֘6d�SߴeeM7`��|��OC{���\m��-��2��I6	'�!	��c�@B���"�а�<�$4l,�!	��c�@Bæ�"�а=�$4lH�!	��ӃR$.k��6,o,q��ƍ�AL��M��R7�1��7�8J�W�@L�R��`��	���Ș�2����R�mC�y%,��JU0�5B&X��zW	�p�A��ƔQ���(�q�w,�[XG)�Ã�`y���8Ji�4���[XG)�ʃ�������`y�4nb�]I�]J��q��(�qky,�;XG)��΃�`y���8Jiܒ�����QJ�v� &X��<�R��1ᮉ�.����q�Ҹ�=�	��=,���̰�=�	��=,���̰�=��,�XG)��B,�XG)�28��&��&,�XG)�(,�XG)�R,��<�R�%%0&X�ay�����#�+���z�*���
��W �U�q�`%VS�L����J*��>�� W�U��TX��R��a=L4XI�5̓T�zXgVRaMs���_�D@��TXM}X��
��+�����R\WVRa5�a�*0�������ǥBK:��l�Nl�\�����]�c�H�y�В-?k�[��BK:��̼Nlu�
-����:��qa*��C�ktb���ThI���b��VǍ�В-�)щ��#S�%Z^�[W�BK:���G�Ƃ�/S�%Z^��[_�BK:���J'�JwĔn���2��ˬ�/S�%Z^�[_�BK:���O'�:�L��thyM�Nlu|�
-����J����2Zҡ�5�:���e*��C�k]ub���ThI�����<����ThI�����VǗ�В-��։��/S�%Z^�[���W��eNǗ9_�BK:��6_'�:�L��th�ƀNlu|�
-��r�����2Zҡ�:���e*��C˵+tb���ThI��kp�����2Zҡ�Z":���e*��C�5Qtb���ThI��k���VǗ�В-רщ��J2��d:����2���ThI��k��VǗ�В-�>҉��/S�%Z��[_�BK:�\�J'�:�L��th���Jl��/S�%Z��[_�BK:�\�L'�:�L��th�V�Nlu|�
-��r�9����2Zҡ��y:�U��T�CǗ_t|�
-��r-C����2Zҡ嚌:���e*��C˵%ub���ThI��kd��6��e*��C˵>ub���ThI��k���VǗ���y�3�U?Q�v�ʉڴs�������=Se��=ٵo��P+{��L�խg���G=S�D�*'j>��u�΋齧6}�+�鿧�V�+s���\L>���\L'��G�᎕s�މ�8�ʀr0��ڥr����r��ۻ^|�k�\L/���p�g��Q��O�x/S٢�.���̼�l�^�Y�6wi�T���Y�Y*�'Pg�<�{�\U�a�dUN6��4Y�zJR],�]n��>��T��KH�;��b:-oh��>��E��,���g�<�R��<�������,)�<�y���ey���.�h�z���Ry���&}�̒Z�|ߙ�1m�(��i��2gD��}�O�L���7�f��e�oB�|�x��6W�|��� 	��
!	��WB�@Bf�B"��|�$d�!	��?B�@Bf�"��|-�$d�!	��ocR$.k��6,o,q���xY���K�(%3^��0��7�8JɌ�b0L�N�$�R2�E",�[XG)����	7��M�ay���8JɌW�0L�<nay�d��&X��<�R2�M,�[XG)��+Ǝ���q�W+�1ᮤ�.����q�W��1���q�W1�1���q�Ẁ1���q�Wi�1���q�W�1ᮉ�.����q��ކ1���q���1���q��N������ ��(%^	c��� ��(%^}c�����ބ�� ��(%^%c��� ��(%^�c�����QJ�
���9,��R���c�b�:.� ��
+���z�Z�
��+���z�R�
��+���zR��
��+��&ߥ�I�H4XI�5̓T�:)� ��+���9�J\' �`%VSO�5�U�q�`%VSO*5�U�q�`%VSO�4�U�q�`%V~&X��8.Zҡ�g�ub�五l���"�E:�K��th�Ys���/Zҡ�g�ub���ThI����׉��S�%Z^à['�BK:��C'�:nL��thyM�Nlu�
-�������2Zҡ�5>:7t|�
-���Z%����2Zҡ�5W:�U�#�tKLǗY_fu|�
-���8����2Zҡ�|:���e*��C�kub���ThI���V��VǗ�В-�Չ��/S�%Z^�[_�BK:��fW��$_�BK:���X'�:�L��thy�Nlu|�
-���Zp��*=������/s:����2Zҡ��:���e*��C�5tb���ThI��k%��VǗ�В-�|Љ��/S�%Z�]�[_�BK:�\�C%�^Ǘ�В-�щ��/S�%Z���[_�BK:�\�E'�:�L��th�F�Nl�V�)-%��e^Ǘy_�BK:�\3H'�:�L��th���Nlu|�
-��r'����2Zҡ�ZT:���e*��C�5�Tbt|�
-��rm0����2Zҡ�g:���e*��C˵�tb���ThI��k���VǗ�В-��Ӊ�R��2:�,������ThI��k��VǗ�В-�dԉ��/S�%Z�-�[_�BK:�\#S%���/S�%Z���[_�BK:�\�T'�:�L��Σ��s��J�3UNԦ���=D�D�*'*o�T9Q+{�ʉ��3UNԣ��r���L�5���:P����S��Ε���S[�Ε���S�Ε���SۄΕ���S�qΕ�`L/>�K�\L/>��\L/>���\L/>����QӋO�x/S٢�.���̼�l�^�Y�6wi�T���Y�Y*�'Pg�<�{�\U�a�dUN6��4Y�zJR],�]n��>��T��KH�;��b:-oh��>��E��,���g�<�R��<�������,)�<�y���ey���.�h�z���Ry���&}�̒Z�|ߙ�1m�(��i��2gD��}�O�?��vs��֫���eq����ƛ���icW���f������kIB�~�&�o/���A��i��|��{%��4��}|��㟥p�W\�Ѵy�vM���S������l��ɺX�BO�~�&`��O�@������4��}�9l���O)4��Xjx�@���������;~�) È0��!�������A����_�"�S@6 � 
����7��ߤy�Zo�]��i���ߛ�	�ݦ�]u�ˏ���E-;%���N�b	3xG!�X���b	3�5R�%�p�EH!�0�]!�X�w}�b	3�5R�%�p�IH!�0�]+i�BdOD��O$P��o�I9 9� IT�a�[R@%@"�k��棔�5�����[�,Ѽٌ7G�X��
'k��;h`��o�J�h�%� `ƛ�R,;�"! S�5�xwZ������f�?.� dj��r3ޡ�r ����f|F@jR�$�\�H�r.�	�@\J@\K �WH�r.l� �WH�r.�� �WH�r.�� �WH�r.�� �Sȧr.�@\�E\��Sȧr.�� �Sȧr.
� �Sȧr.6�� ȧ�O�\��ȧ�O�\���݅��ȧ�O��@�ȧ�O����ȧ9 ��5xA-��Os@>�j�_;Yd��W����G`>SOR�� �����ԓ��8=H��|�3��PN?,���� �oR�Jx�X>��8~�JS�����/���T��/���|�����A��#0��'špz��a��g�I(�$~X>����	4ځ�		M�s�cw!p��!�6"�v"`BB�C������Є� 0:�hG&$4!?���!ڕ�		M�^�c�v&`BB�C����	��Є��;:�h�&$4!?���!ڥ�		M�k���>LHhB^耎!ڧ�		Mȫ2�1��1��2A���)�S���&��/��}
��Є�tC�O����c��)`BB�)t�>LHhB^!ڧ�		M�K��1D�0!�	y����O����c��)`BB�zFt�>LHhB^���!��.��]h���>š}
��Є�C�O����c��)`BB��ct�>LHhB^7��!ڧ�		M�k��1D�0!�	y�:8��S���&����}
��Є\' C�O��k�c��)`BBr}t�+Q�KQ�>ţ}�G�0!�	�.:�h�&$4!��@��S���&�z$��}
��Є\KC�O�����c�>LHhB�a��!ڧ�		M��w�1D�0!�	�v:�h�&$4!�=B��S���&�M��W�×ͣ}J@����)`BBr�,t�>LHhB��!ڧ�		M�5��1D�0!�	��8�9ڧ�		Mȵ��1D�0!�	��:�h�&��g�9�q8w�Ma�IM���'�Ugo[���?���}|��r�
�3�O*��l?�:�������%���9��m����N�W�+0��;W@��܊l���_���K��S�t���Ui���Y5W@�m��D��v[{���=i��G������:݊�^��E]�YB�yW�,���m��̦t�cӏ��K?����Y���t��ڰl�*'�yk��t=%�.�.�ya;���?r�!���3��$��eV�h2ɚ�h�.>:�;������/��*��ʒ��S�gM]��Kj������j�ߤ@�2K:!�}g�ƴ!����-+����3ۏ���bq�n���I��7N?�g��|��4�3M����ʣ�@��xC�2����ćK|0��ćO܀�Ű�������[Xna�Ű���[8n�R����g������9���ajpNw{�I��9}�᧜��5H_���}�㎿�:��d&9<5
{��Y�N�HB$ڠt��s
d%@��I��a�@�г��M��D^"�"KG���_�v�Ν�"�BF���^F�şw�U��W��a�]ܽ�L��[4}�޽e�o�����-������
ӷ�r����z/�u���V7;��Y��]m�?ooc]�PX��:}d�ַE�Z[��#}-ٲO_��s���%�M��4�C=��4}�p��{����]��>/��n��v��È��z�pI!��mW�ӹ����o~�b�Ssu����IBo׫��H�y�����뤻�웫��޼�ۿ�nV˫��m���j���.q���}��Mc��v����G��nW��$�\onV��&�ᵫ�6\x_��+E��I�Ҕ�[o\V�`�6�6��K�^)B�=��/��K���t�HӤ]�nG��&K��v�T��p1��v�m��ݷ����"T��E:����/}�����������+���|�壂}{���a��Q�=�@w'5}�>$>q�x���Bq�S���_�j�;��3��Q9��s�
I��;yy��X�2}�X��-O�?̖g��S�����:������nu��I�:~ؤc?l�Y��*N3�'Z���4���7W]�^||3��7��7����]������b���+SR��uy��.,��-m�T�m[떾	�����Mʵܽ��flkʲm�f�Y��mZ�� 볔���cK�Ж?�]컪����Hf����Ц����gjڛ/�Y_����!���3�1<�E�-�>�;�Cޕ}5���7�?E��6����4&_�[]u�XD	�(҈ڧQ�vm�j��L,�m��\̓P|�l�����q��R4E�Cj�u!�q�YfKkB�l��]M�Q��js�i�Lݦ-�<��<�iX.�M��]�ː�e��;���|ݬ���x�J�5�(�O���zP�{��i{y������s/���f��m�m����{�.�§��_]�#����N���Q�	56+��� ��Zv�m�UYKM���`y���WY�&u�HY�QF./Ҝ�S�ұ��H�<��l����mV�y��"o�3���<��\TK�,:�]�>>}�Y^�Ͳi*J���֎�|��i��^�������닏oެ_���o^��{���v;��~�.n�ŋ����v�b��������?������f�>"��ױ����}����x���e�O�b1f����Ù�}���`T�����v?�n���˼fA/�K�z�t~����(����a�p�l����5|�Id|���m�p޿���{0Ϥ4�7EGY�B�u�Y�t>���|*׸�Y�̳�j�3����&SM2��ؚ�-������4"Z��N��(�Wf|1���z9��+���<u���4
�Vz�f�[������U����Ư���K��e^�7|���7R��9c���v������H.�-O���ӰI]���J��}���}�*�ӮXgyirYrW<�z��["ƞZ�/}�ܽ�t�żL#�ˌkC櫘�*��d�뗑����;�J�s#f���99�`JG�:/�y?�?ś�x�{?�ns�]���d�/?k̗_�����c�1�����O��������x��rV���W��?o����&w��{���������\�7r3\dO�+�d^�������g���5_�9�Ӟd��n�/�������Ҽ��Q��c�(@��p�����M�?��@aS�H�y�7�W�c���N�O#Oن��Yw=θLbG���w�g���G�d�S��i.�mY���/<�y2є�_Y��*���pgtલs�r�{����/����.����%����hs��9�T�0��c�q ��a����ki$|Y�4����a֘����ȟZ��������]��r��6�v��e?�{�.�n���V������I����IQ��^��w�Nt_q������{��ֶ��Ó|���2K���Y�g��a�7���U�{7�%��f�� ��_�?��~��5��þX?�!�G���9v�pyl�Q�O|����S�_;KS���b-����b-��DW���*�����ÙG=�<����ۆ�y��u��V*pW�b�f�ã��?�U>h|�Q�����P�n�yԹݮ�c0��
\�����wEm���vf�;�C�v��]=�=l�+7��s4cB�*�F��8��NS�����T8�5�����:w��ڸ�Yp�l;K�v�l��[��~��NZ��� Cn�Q�v���\��,;dwQ���<s(z�|yVw	��a��:�]�"�������f���ׇ�t3�c�����Y�6W_m�����V���ˮ������w�ݮ��p,>�PK   J��X�J �i P /   images/43ea4950-057c-4494-9498-aa922855ac7b.png *@տ�PNG

   IHDR   �  �   �$   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^���e�q�	�u��z�M�n��4� 
;Z��ӎ��w$�ҎF�!5����5II�FԌF+CI�4R� 	C�h����.�e���{���8q�y�^ջ�]� ADU�sn���Ȉ���<y�I߅��w��]�.|�߅�x(d�o[�v�#gϞ)��%� P2;Z&����/��y��k�q9;�����y���ى`O�� �ᜎ�BZ_�G�Z�g �7Н�Nօb+��;��t`&#=Î�����(`P�p�����j�++�]�b�ĽG�ΖRiR�G��r��)w��Nэ��.t��b���#A��n�r�E;��N��h2;�\�,��&�(ǎ��c�����o��R�C����N���RA�BQ<v��[GEeQ�!�@*�\���/�b�5�:�<;��նv��muş��Rb�THM5��ju���Z���#�����oZ�\��o;��2�������F��F���N�yk!tSgZ��*KE(J�J(
('���2h���l�~�?H1[~� �4�7i����F�������?����(����28]/�O�,`t=��z���Y����RjwZr��o��R�\8Q,��Q.��y���ψv�I~����V��6vf�̡������'��P��]����-��򚒰;~o��h;�V:�=������o�ns[�.�]����4;m�}�t�ِ'^n����T�_���݅��'fg�,Z�o��[����M�Z�O�;�OH�7hH���V���!�R4��1r].�oCB^������5�n�}�z��y�m�:4����Gݔ�E��:�3F�mu�W5F|�T.���������v�� .���۵n�ժ��n}���w�RH����wO��1�>h|=���]m��'~_����������߫'��)��k�����e�����|�4:�ϧ��~�޽��C�t�''ΝK�6����j5>��堧�w�p����߃J ����^��
��zԑ�k�:H��7�H�7�<��t�e�i�5m�#@�h�žʣ	
����GFGijj��8빾u�ӈuU@�,-o�7��n}L�2���`�<����b|g����KѹԵ<��;��y"l��nw��l�ssc��U����p�.~�[b|���ex�0�	�4ó: \�y�\���3��iyd8��vy�Oy�瑾�����0�?��FZ 0�6���L<�J4$5��fЙ�tZ�V�^_�QeY=��A_�o���.T���7k����v	m,/t�Ȓ���S<P�S���f`¾�`�� ol�c�Y&�'Ǹm�.v-O;?��q�r��A�1�3ZŒ�gS�>A�NP,U^,�K�����x�ȑ��[ �� �UΝ;wg�Y��Z�^ocC�+�����}o6�0h$�|��B���Ac����(�;����y���,VG&���|��Nc"֧���#.����luS��iubb�禦��=x��fV����媀f�{������wI�s���Oao�Ȇ1j�v�+̧Ű�-��e!��6�)[����������uأq�6:nM7Ϧ�m�ua�����B�8��V�q{���=�Ri�U�-�7��$��n�yS����~�����F�6[� �LJ1D<�y;��(M�R�y�\J�P]��H�m�nKu�,�����R*�E��T�RɎ �A�R}]�!C]ku�J���X���V���;gʈg.�Hŧ��+�_I��Ie;�g�v�B��B?�pvOg7��w����g2"rA����T;�v^�5�s;��J�;��G�K��9sf���}O}�A����յ�J��G$�C6ܪg���a	�{C��4!�|�'�b��X��>l��P.O���Pl�R�߭���R�O�|��j�i�Z�6;g��s�RqI�6�FƸW<�)d��w��wJ�)�ʨ�!�,D0C�7�]�d ��|�whH�-�˝	$Ҩ/���J�#���n��������-�����J�Ǝ�?��{���OJ��፶�M�)"P��ƷU�}�*|L��*�2g��t���_Hj�e����f�ͬ7��Y�ח��T,��)czd�\yn�R:7R��(���Z��rY��z���ڬ��j����v��2�I:Y9361T�`d���x�:$i����v�O��c��A#F��W*=<1;�w���~naaa5�����\]XZZ��ը��V��#���͆�é �9�p���u^h|���tYC�	5+�7lһ"�E���y'�G|vXo5��??R�|�T���x�陙�ř��F�p�7�UVD���9ӜY_o^S]__�Q���n]�])��ʒ�
1���9�'�/��o�$����9���%����yytb��/���{��L����&��<yr�R)���h��N��>	ܼ�����BA珄8y!����u���b��D�t$��]�(��a����_����]?s9�A�/�}��=K���77�?��OƷO���np�ǧ���q�o����Q �`�����������,�*c���M��������[�2_u�7W	&&J�����v۷�p�Ƃ&|I1o�p0����c�dF7�~a�Njh���ȣavU�o��O�o��ׁ^��e)�����{����Iџ���D=ah � �����y�������As��9�N��F��}��s�,���j|���|�f��W���oL2��ыuёs	%����B�SR�Fa\�c�7Qy���}!*?ld���j��ybjr�_��-|n��׷�c~����cӏ�OL��8X�7�'��e��Ч���Ʊ��-�v�Q���a�0\v��;W�P#�~K��u�&'����3[�o�c�Z�my��y����U5�����f���-Rl%�|^���P�`���vy�Z�<�۱�Jf�B��q�.���kf�KW�����/OLL?R.>�Iș0�>?}���,\����,:���v��ٟm���#�j�}����,��U3��������;��G?����Rq b��+ �g��=a^��]�f�Y9��!ʄ�Co`�Q]j���N�N����ïf��>|��b��h��x���)�p�>�����ImD�	�PF�ǎ�X��f����w��g����V���μk;�j�v�7��woV�tߠu�����HpL��Y�*E��cC(�סּۥ��,7X7�Z�&ٷ_��������K��gWD�9==v�R�|��n/R/��{�<OW��K��c�,��~]�^}�J��.�W��������Ɲ��y�k�oih������6)4_�	(0�>*�iZ:y)�0��;�K�f���U*�o��=w���y���p�P��&����C�)\^	����c�hy�q��ah��>F�AD ��P��B�V��������Kcv�*�U1�J�{���|���^�g������b@>-�����>��@�{䍪�r����[b(���F�N��Ӫ�?ֆ����6�c��>o���SȂ��)�� 7�W�޿xr�{�+n|l�j�[�(6y���=j��p��5�B1J&e�H���d?{�=K��#4�F��t�����+�s���
H����,+�Ո����6�7�|p�"OX�����f���94l�U.}��4���2b�Ni����Bc���Zm�M��q+v����Z�v74�OJ���@��r�H��<Ƶ�֎�/��Ǽ��w��B��_.�6b�*�J0U���˥u]������|�L�a�5/�' �y��������FY���k�+^>]ޗ�*pE�osss_��|W�Y���jL�07 G0�Y���ѓ]8x\( G�ؚ��Vc�o0=�����o4��N�PCW:c�b��*�b|�o^�ls��ہ��(`xH�6����呌����|�ˆS�}ǚ(�BN�Č� ��Uݬ~hcs�ƫ�]1�RG�����V��V�y;S�{�h(�b�7� ϽA�?���B��|����s,�Td	�R�[�W�me�
�v$(���l���8�/���]��!�A �zB���y�P��k�T��x��b媭�]1�///�����ݡ6�橁�t�e|�8�]��	A��-�����	0�����e3[!���&ʈ�[�FxR�(Ք��R�eyn���0Z(w���G�������T��.���.�L�aP��E|�'���s�{F��M�(��2�`/Dl�#�9s��sζ1������F+aj�����/+�;vub�+b|¸��Mb�����t��{)���e����\�q�n�[��ZGD�c(��^�G>�+�JJ��½k��j^��@�ژU�Z�i���V4:x��m ���o�\ۤg�/v�4��]X##q3��-��h��Qk��T�k�0\�[YY�߬7��m�ޤ�4���	T��@~Q��0��(�9z����øó�X�������B�ߙF�%uy��f����f�֯�<At+�k+��u�B��ݞ����Ӂ��0Ѿ����Qli:�l�݊EvO�5IJNC9�:�S��6���z��=k�|O����u[`bqS��������З�у��y��"���7*h�!���,-C3�1d���|=�3�nwn�7������9�+�ν���^�>�R{���cZ��m`K���q�JA�U4�ͧe#r�d�sy��-Ս��.���{��W_]=� �����C�+�'fb�j�K�p��4�g�!��2�Y�S���JӱG��	u�㉰�gw�{�x�a2^P<o)�n�@U~Om��޵��(��ID��x��M�z��bi�vg��JI�'{�)��Y(�o��j��r�@_2��7$j�#�|��n?��:=��2�HF���/��U��د��fm�MW�Y��%�n��T��x����X�G��y������<xZ�@�4�n��(J�-�.���Q�փ�s=��|��\������Nx���+������]Y^��f�6�	#-Fud���b����Ӡ��0�0��Ҝ��߲;����ʍF�͍��\�'�^���[��ʋ���{o �kMy��Qލ�zz@���E۽%����+h��t�x����V�ul�j׬�����ųZ[;uEn-;�̡��^��V���r����ldC���ډ!�1J�>�e�	-�@^_��.���l�@FŘ�B��!�!'Յ�8�:�&��oT?���y������l|��:�M�!�����v���)q�_�����~���m�$� ����
�}^HC�\G��V/k����,���gO/~h}}�u��;v�����]���aq}m�R.�h#u!x��
�q1ȷg{���˧��r���ѕ{E���ʹ�T^�����l�o��o~�ө �J�k6>)�<�����%<�z���|$L�Jc�0B@�\�(��?��`��t䶇�s�z�.�=���ut��e�RaD�UI��g/75>*%� Q�z�H��F+�V�u���s�������Go���>gn .z��go=w�ğZ[Y�����m�g�Ր��&<��\`�!"�C.`�� �?3Ҹ��=ϫ6��f�$Q��Y_%��0��[�̮Z��յwhbvE�����L:��U,��z�mD�Ʒ���'����	�!��=>n�D�]�0�	ф00<ش�UR�z�B(�?����YqM�,@�/4�.������5�B�o{J�������s�_������S��SS��T�!�^�@��Ley�前��޵͵[�7��okkk�[��K�گ�׆w<-!	i[:ں���_��?��v���10��䤿!�8@�{�/��3X��Y=�\3��Uetlujj�w�w�����+��ڌ�5_&��-޾����n��'���b:d�ftH����z�r��X�`F�-� 	���AB��a�J �i�}�S���ə������dQ�V6~Z���}�r�bˣ̥����������FǾ11>��he���{��)6��F���V���l�V�v����F�~W�ݺ^C�.4oW������k#e�'ۅ�v3��S���m�c�C;x�B\�ne��r09g�ށ��$�]���|�#���{Q���g$��M<7?��s���y�u�d�B�w 1>%��)�o�V�m2�"�����g�ʌO?�FΪ�yB�0>��!� +�?���a|:?��2���ax^�+�s3@y6;�.�,?�e�7o.@�q�^��G�ľ�b��2:2�Z*�7��b��jj�,��
i������f��¤h�b��z��������Ė��:1�P<�ubǞf��:����h!O ��h8�|LȀ���o�lD��U*�:J�������Ѩ��������]��P�-߸���o�Ɵk7�{-h���iΆ[Ʌ��oٹ�,��	��근���ڤB׹�ke`���:�Q��N�3:T0�g�'ۭ���/���<%��f&/���@�GЪ�<@�(ó���%��:�kf��lW�"u����O`|�#Dq޽^ o|�?��AA�Xݙ�CZތ_�� h�o�F�娺��8w&7zh�<J h򜚞}ezz��.,�sss/X�� }n� 1;��|�=�Z��;��4kՒݧdX����P��
�<ݮ�w&SDN#f����P��r���ȉFI)��bb���j�53F����C^I�)So�8�CHiQ6�s�p~l)G��0B�#Bh5u��W��Ŏ�̮ѣ9����|�Fm�	�d�����eс�7�4~���(/������� �fm����ع���:����B�+��!u�������c{�������ggff^��r|	��8{`uU���Q1{�����1��7����y�h�ݓ4Ad����<�� p�C�а!���f�\_Nk�,�b�c�%��������&ifz.�OM��I�6��[��ѧ&�-ؚ��!
��*kvnl-�'itr*M�L+8��������༩�d}e5U7�Ec�h�*?���Z�,e�<irr�Bx�v��r�ae���8nɃ���kvn��a��c��ח��F�Ά}���o�ͫ�v}ff~����3��Ѥ˂>7C��ҙ�7�k��n}B��4[�i�5LB����[� �^��t���ɸ�[��@��ѫ}��D�ܮ�\�;R���sieiI�����R�3���-�KD�g/(UCE��`ZXX0Z�j1�n���tӱ�G���J�X]S� �V��T�њsRm*צ]2�م�iρ�ifnV��p]��]�P��L��ϦWO�P�Y3ZS2,���ƻ�%9)�26����g�l�=e`�D�����auY�:��gymv�J����2�`'�v���f��F���y�r�^x{��s��4�����ߖ9��F�,�`TǸni�AZ��c�*�T��V.8D	9: �nuc-�;}&�d���b
T�F�a��I߻o��iy������q���RZY^J���ehM[���7ާӔ��>���B�����;����m��-X�d4�[�71d<�����Eձ�
,�([���GY{��7�v�8�c��Q�v�yI6�j>'Yy�	#�a���Ǽ� �%?���N����L��eet�jw[j�3������s�aH�Q�4��MM�ݛ���n���P9��x)���5��f��#��Q���K����WFd`��s���|*JW <6*E�Ɩ�����Vd4�k�7օ����i�W<k�R�a�x����(1�.�ڈN f���Z-5��T߬���bm��C3Y�Ic�1k׈�7b�0^���F	�:��+!l�X����# K�����q�1��M����?��ˬ��3�Q���.�H�cv,if�L@[�S���Ïdø|Dq��M.�!ah�k�Z���Q%�4�ʌ,o�q�kQ�G�� �qY>Ԏ*k׳:��S��и��uks}5m�&k+2>����e|�:߬*6�0Ȍ��=��XQS.z�@���e\Ķ5�UOX�������F�}&[�FC�*24h�T�Ԍ�թs�_�Mʯ�s��?xT�a(^�XI��f��6�mx�Q:$E.������2"�:�����~��)��f�7�J2(M�z�N�,�8z�(�Q�mܭN~�����2��I	v�*1�
H J�I����Z�:e�.-�:º�(�6(�٬k�Ï�R�Y��ڴWS�����s��"c��ȸ�4�K�Dd�A�k6����U�uT]>T/)����Q���bTT�q$`m���:v�͌����9��:˦&%��ֆ��Q�<�u�N�����;��j�>�������T���t�d����J��y��T騼͔zm�f>6�P�lk����A�sa�df����\GK��fQ;1�դ��c���T6_�dx��WF����LPx��o����غ]�ƀd8�����<@(+�M���#�F^�_�)3ȶ��N�n�)�g��s�j���ڑSe��C�#/�p��x���E�X;g��7ƥ�ɦpn�y� 3�R'}�:�z��P�'�~qTL��+G�`� 3S�c���ye�hd���q�^���#��{�f$�p(�(��0U7^J�D�m*A�0�x$�Σm��r�W�����7�ɳ��U��b�y[�?ꉶs��"��6b���ݼ��)��s��0~��S\7YQo$m;��kypc۞��hK�Kj�E9���6��FC��\(��Tׄ*,T��<�	��[a	�2�TF�y/���2��Hv�N4��&�	Qv9��3�ҳ1>� ���dƆ��nfX����~@</ƠsLc��}c��� ���͹���E���f��N�w��m!_�2b�:4D�n�C~�F �+���Ґs�Ax9�G̜Id��� t	��%���C?盫�Pj�;{���H�zi�h�<�Z^_Iy��PfK�*I{#*4�����}Z�9eLA��$pL4�c��U3���u��\�k�e�Pą�A 墍����xf�s��]wT]v�E���P*h���4b�4�r͟��bЯ{+��DZ�j�o9�¬��GC�h�Th�g�P���H�-�'ы%6C�h�EJG�Ub�� @}[�i�aP���RZ>�h�3���E�C�R��s����%�o�5��RG�{5=�^��"^��-f����bG�s[��\�'��~���-&�H5Ѓg�<K�����נS�L痜w�ĵ3gΤ�bJ�Eu���6=yP���ty+���L^qD��Qv��v��>0��zQ����5�Q��ꊈ_�	`(0�t����;ߣByT��ht`,Ap�Z��W_}5=z4�8q����ϧS�N��"3F�P*0�|�<�X�.Z�x�Cѭ�q�ܹ���W�/��^y�t��1�=�N�:��?�������mkr��^Q�!�Y�Ǆ��h�WϝM�?�Bz�ӓO>�>��s���^NϽ�bz��ұ�'y<���L�Zg�?�c�� ��ρ�~��u�,TTW��`X���)H6����.3��p�S�J�Ӊ�p�����7ձ�����Ԍ��V�ZO�k������aX���f3mn�F�٣�-�166f� �ESã�`��s�B/���F�W�ܬ���ʹ���6�{��h�1�MVx�M�Q���%(��V�H�u&/LdTuG\��i}C�ա�75�CD��@���k}�D=�A�x������c.�va�E`X�c��f1/�p�0��y`]� �!X��-�f�X ���pH=��؄�q2U�Ħ�"^:�K�77�0��53EWk�E��Qgy����X�
-4V�p��dȵ6ґ��v7C��3y4^�����X�5�+#i|j*���b8ޓ�ԐYV[*��i|b&MMϤ���!��!��bx� dC=юa ��"=�c44��B�ex�¤�Wh+��[��8R��q�x^`2�#��
�a)��q�FBB�e���7M�3��ܖbl4��L((��X�A�r�A3b .4����ǾP�o���f�y�����PA<�ٷ=_"4�W�a������Q_�&f����l���U�Q�W��#��z�i��-�JO�L�,4�ę���%������v�2����<�$+K��\m	�:��r��C�b�15|�N�/4���3�7��,p��
�{���A����w���C���o 8���ѣ�5\.�0Ɛj�+�c�ME�(����2�C�[Yqst�4y:�s����!��ȍVӼbm^F+
�~���L'N�1O8!#���5�����1hv�q�Ao;9�u ����� MG����f�`t���$f���ƞR�3ߐ`&�*/oh`��FG�2d���sҸ�Cb+�.
�׹O����}2��4>6�x��^x����O� ϩ�9��փ}��FZ��0�;�E�����M���]Q�b��Ȉxq;y1؏�O�UņO>�L���4�x!U�NMΥ��y3p6W`��O���/-AϮ�|2=������A�fV�V]��z>)�ohL�����4�3��Ȳ4��`^���!��D�`��Ɇv�Z�ǲ�?��hT��(e�iU��W��HO<���Ǖ��1a�,�")�	��s�d��C*�XJu��C�{�1�*ڵ���E��zx��?��;)j#�I��N�S��W�7y$=����F5�d�<ܬ�A��M�IB6�*�f�m0�bh���� �o��}�N���o�Q�tt#1�f�D�%�a���#�_{z�s�%�^`�6�vz�g���9V��jL �*'gf���]ilz*UۍN��^G���;��r��ַܙ�ւ|�֮h��̲A�e�k������������`fn����6��W}�J��!���`�m�s��U��"o��;cZ��Ď�1��{מ=��׊��Ç�I�H���B�	�E�H̘�ك��e6��{l�kFo�P��j�ntջ������O��_�4@sGX__���j���L��
l1,�����6�z�%�~���Zh9��G���NR���6d$�.�X߰�Ilxc3ժu�.���o���k�^���1sdd����Lyږ�Χ�gN�v'���
����w����܀߳����0��d(~�.�bk��s�geq��!YP��g޿�Ś�v�2�ȓ����oj;�	/��d!H�`P�
!Wxw�K�� �1r L����������*^�؅���%@�w��o	?���Ӆ�7����p�4*��%�����9#��Q^�0~�������J�(3�&�D�-�H>��E#>k�,����þ�-u��#�9�uy� ��1T�����4<�=��b,�0�n��'����g��Q ��B��� 9���30�jy�s �T���F�y�L�[`@�ޞ������s��2��U�fX-d�p���p!^
zy�y�lW��43	��^��o���*+e�����es�-QpΌ��,w���1��⋶o"�a��<����l����9-����3n��U�i��� ��=�aܜ�?�KCiC/�7��v�(>"dw5i� �v@�q��z��F��>C;���OM
��-�0�A��y�C��� �9��~�T˥���5�#/��BYS��¬sd��P��-Բ�Gh+�(�{�d++��e�2����Թ<���Q��=�Ƀ��F���t*�'�$dy_}T�.!��ѼN�9�j�-�ӹ4���Fڬ1�����+ă���N�G�nb>���G04���?y^�\���������	;���]���P�0�; �!�{Xo�ֺ�b�P���`<R$��rk���d�w!�]"~
����^ݢc��xTiʶq�(��0����8��1KF׎ޡ����e�z�H'��4��������3�v�MT �҇�ȟ�{= �<��^\��!<F^lЋ��@��1�u����D��9*-�,��˖.b�<���,�n�)�ØFku���?a�^:�ڳ��^�[kB�ed��H��"�.ވK>�_AC����O��,�#����uJ�Q�l�[6�aF�R�v�eBN�{�8� �.�5a������0��2��Az���~�� �l���p�6���@�s %��gO,�qh"M�o5�	^&��J�Ly����Ϣ�3'��`��y�Ǎ��X��3�+3f��mB�4 ��7�����lA��.h�!�Y�z�s��lW&�y�o���m�;��d������B(�By�� 7F�>p-SNV>� y���(�c!U� ����:��ZC�{,5S����2e?���2��*>�;���CRr�c<�x�(��QO��om񙕅N�:�@�|�]�ߞ�i�-6�T��]V����x���i�6ႜG�9�����͑:�	�,Ă�� �P`U� .�,o�1�P@�y�x1 ����y%�-u�fgm�\`f�4�Xr`<�P��C3�Dd�Ύ�	���)ʕò�v���6p�t /��q)Z@\�:F��|`���?N@/8c|����N�	!Ȝ���y�4��ը��(E�b]��Z���X��v��G�f��F8�E������-گ'��j��<�o���G:��]��O[䴳��H���n�:����^�V0�dG��z{����N�ٓ\����!���Zlk>�,^�1>Ջ���c�_�!q�2���8X.����i�hC(s��s��ᅿs����\�c��|y9_dΰ�RO������I�0���G��s�N[h|g��Г�hF�c��A�S��% �/��z�;��_`���vg�_l��Ł`Rule ��`z/���a�\���h���۹b���G�1h��f�Wh����X��Y�~��Ӷ�,U�1ڑ��"���P1fQs�K)�'C��Z����a��2D�����|	Æ�(��L��t�"?
����Ʈʃq���{"m�1;�XF�� ��9��[�;���2^������ v/	�
�]B�y����1#4P�&������8�|M��i�R��,���mk��<��8J
�	ڑ2�A�J��1�n�wų������Yn1�A��V��73l��BB��f/HŔ��?R�߂3œw8��������,�x>�������q};��-�O�ݣc��giԾ�����(�Wʻ�.N���2�k���>)bel�L��#�P��^A�0~��3����~�A��!��H��z}L�ӧM9)��-:f�7�<��qn�ˌ�3ڙ�Q���� �^��>U|���B�>��t��)�it�`�s���0zB@�6��������~���Z�i�@���y8��Q6ʓi y,_fx�?��~y||��OLL��ʭ؅�K_h����b�I0Ø�J`�kX*��� �w�#��P8�$E�(����]&~��H�F�z�d�0�M���f��˒��o�7H?���6�ijC���J�*�����+�'G��ky��H�R��A��a��u9Q�D�i�c��o&#;������W��!4�����İ�->^f�G��:z����,@.*g|��ܲɴ�3�9������n�B��z�*�PÈ=s+�(F+�Y3E���L�ƣ��d�c�+�b�҈��.V�u�t�u<�	�=O|����J*��~�ƀ�F����m(����kUD���9ڱT��Q�����1�^o+F�^Ӧ��T[
��=収���zb�;�mci����kw�`��xؼ,z�7��?o@��J%��=m�#��t�mk��e��F蚧�q��M���M�Uݒ9��]@d�N�`k�6�R�[��Ꞓ��S�N��Gn�n@67MG扅��/��������o�'>�# �KBf|w5��ow��˲$(	������4Rm}5�y�D�X[��ǳ]��0�Ch����4�]Hcxl?t�1fÏmQb��0��>݆�a����|.�>y,�o,����ߴ�Ù�߄��s��5Gn��FR���k�h�ІP��Ǳ2RJ�K�j�i[�9"�fE���(�z�����k����q��� <
I>���n*�ȇm���zZ�œ(^ސ�p����c|������쮆6iKe{������U�_S=m���e�7V.��2a�ᙡgzm�-�a�8󛇮X����[~�~fu^�F9`ss�O$�O���Es�aw���׫��h�ޭ�ev���&�S�h5������JQ'�7�6��a��)�.�Y���TUY�F�P�f����=������CG�7�Q���k��Ui⨑
QVK�����ڽ����GG�He�~����R$�����L�z�{��Ԃ�D�xS�����c��iXy�GD�����m����H�}��Y6�y����o�-WͶB�E����0���_��_O�<����`R4&1 ��NOO�����ZH�^Sڷ������5d�q�VdKy�r�̩t��+v��m&ބ� ��&�H333��N�>mݯ���Ca$�A��ɉt��a�;MN̦)�����>I��V���]�?599���k�*��/?�S?U�tը�7���:1��z5�]O�͵�t�����x`T^������ �^��G���$��R4�M{� /U�����ܼ�0l�ޛ�#�A�ۜx/�y��������_z�_
������M����b#����C��n�9MH�қ��s�(<�$M^R��/<�\z��o�SǏ���m�	���߾���v�?t0�ٳϼD�Z��Y' ݳ"��u�W^~!��ܳi��Y���bH^p�fƲ�v��g6���ڕfg�T���t.��75�^Y:/~ys�Q�4g��ޗ���ɸ��d���tp������O�^xN�H��-�E���L����Y�t�_ `ʪm���C~idd�������:;���Km,���Z�ga|����Q1,I*"H�%�K����g���89� �N���7���˰x����m��O^�(C�b�F�� Ęy�:��
���-|cI��XYU8���e�uu�����`l���O����Ĳ�;���Q�G��2���5D�w��wGT7w)��Bǥ0�<.v�� ];�&U��A^�lɆج�����##�t�Q���a`�1���^{��ґ�}�C�e���Y�[�8W�Ļ�ժ����ұ���΍�űl�#ȉ��[޺��x.�WY�}7��k��K,؂�N��i��!`�X#�αUb�lKë�:/�m�!/l����O��̮ի�u{.�W��	�k_�A�����`9G���0y},o�o�Nm}��omy�f���J�Ge���(և]&�M
�Ƕ#����tB�F]4l�Đ��w\�a10�{�y:�����F��몍#����N c�ónVW�{7坬�+=h��t������A&S�G>�YF���q+��L�u��WΧQy��	����!n+���,��.�����fx���$U0>�lΆ����0O�j�a4Tq��,aK�o	-(Ή� ���J���U�l�%�X%o�8�Yg�*ob�&^װ�˻ו��0x��Bz4��5��L<iÁf�-)��^������R�lQ|�o�����>06k����ӣ�.!���MLo����x&4�FR!��G��Fψ���Y@�^�H�t0�C���*�w����+�dE��Ͼ�.ީ���`����D�z�̫���a\�M�tF'���TW�bۊ�%���u�5�ؖ��쾦�ӡ�hy����\c|��L�B�K��0HG�:X&�1$����ļ�lR
��;���W��r�)�ճ���ƺ��<�Ϭl��D��3���1�]�(h9=@Y���0�8@}>k�%�w�M1D�L��B��JX3ӭu��7���S�1,uʈA��ĸy�s��Oi�#7�:�`�kJ7��yAA�bDaF%�l�Plrg��9H���My=��Pxՠ+�k�0��axm5�k������RA�x~�R�).8�ݾ�������!$j5��m�#��}c(�	�fM�R ��G2�jL�>ܡ8f{����!��cQLgy-M @�L��� KI�u�G�<�S��a�saJ����[���v8�%!�`O�1�7����@I�N��)K���ꏷ40�b)��xHx��h���e���G ����o�,���J����Q�B�����}�@�l-f|�&:+ț��[�i@�r�H��5̫�5�U��I�Q�z��g�#�Q<� F(�4�%��1��f��j*ySTA��8�e��Y��)�L�|?�^f���8�7FP'��@��c�%����%�:%K��G*� �`و&B��&�y̒#/��U���p�I�+m��yC�k`cR��P��X��W�B�ht�y���8�,��<C��O�p�3ibBǩ�ĳ(�M�?��W��d�͌٨kO浱
߹����m�:����(��<���,÷Hl�L<�9Ő��i��\�����_Q�D���`Җ���P\�"18�,,���!jL,��
��ձ d��3�k1U�m)�*��A6�]zM����@��Y����x^}����*OY��93���9�ߐAVu�۪��&Ƨ��Ht� ������0�2��=�2�o��j{���3���湳�|T�[dYL��Â�@zC���T�A�uC%���4bO��]��ԓu<Ot�����B��X'Q]<!gu��[k�W�U,�ʖT?hz�Y[+�6J���#Z��5�������|n����3��t��@#���K5���z����ц��?��F阬���r���sijvO���L�J�LS3�Ҿ��5�_���?(Τi��v�@ޓ0<ll*p֐��'�k�����E��Q_�i��(ՋgAx�I�0�s5���h}���z��g�WkH�rE�q�a���a �B�>�3���4V�rݣ�j��@�W�L��m3��{`�jO��>Ft:Xc�@{EӼ�=R1��S{bMu�IRt\nb��o��0̪����#��3b�<j���NJ)�4��C�1y.F���xnZ���p�~B��4[���zR_Y;���v��U��/����]J���8fm,G0KjJ��?D�6Ӈ0<�(�h֬P@:n�z�p��klX��"�5	��0<��ȫi_y�E���CwTJ��{yk�F�|��7�뮻�h7Z�[�q@��a����N�L�N��١��� �;Z�1X�q�c��}i��}�p5ȼ6��q#���y�9q"��,�����I�x�����T���,��J�6�|/�o��3U�O�8�IǪ�В�I�L&�$���u2���W��}IG�q�/��'�5a�ǢРc2A�B�'v��[ss���\�w��)��m_��q��D�.6e\.T�isؾ/��32���?��^ B���xV�Co���Zסw x���v`�</��f�2(=���0:��H1Rt���Y���h�}�p��+�)�7�2����cyܟ�����E�hʒ1#l�Q��-�jU��d�~����u��f�	�8��o1��g�+3�o�g�S���d��=ax���e��E8���*�9p��0�Hc������ ����2�w-�����n����a���J�"�i�^}+��*lr��Q�X���3�C3�������
�'r�~���#�ȇ�D��.p	܃�m9"@�& ��k��2=�k�c}��)�� �yt^P:G<%^ή���6����ЀS�dXf �gF$:����'U��[��آ�:������Ɔ�drA�ȀO�[[um�~�Ui2G��`�UQ�� ��g|kU2m�6Ӊo�4 #�.�b{vI��:f������m��g�g�~jff7�7Ԯ���%AO��E��Pգ���=?�lB�=uL"�ًB��l(qrݼ�b�I�C�M5��G�(��g#1���T�ZkG�� ��B	�":(��# .�\V.c &u�� W�{�� 4�f/_�ۥ8f��ԭ�5S/B\İ� �`=ۚ�<|�K ۥL�xE��xL�m=��B�����M�5�^�.���LHF�7&B�,;<��_rVe�Mۡ�<���)��D�̣z=��<:v�����h�Gɫ##J,���#N�v0Tf�RLc��s�ȑ����Y)����(�p���m�D04�BF�2�'gBs�3,0���J${ =C��pK�(o��K#0O܆��Wf�pʰ^��D����J��ϕ�9�1X�s�\�m�s��j(>PFe\���R9h'��Q`�i���+�j�b��O�#Oې�+��ݒ�u
��DId��x�᲍���u��h�)ş& �(:���E���3����@�E��r!s>ˊ�p/�3nC�!V�.! I�ڦj͉�ͷ.<0ܪ��&�#�F�Y(V��j�
��N ��bQ6�1�͊��Sk<�3����|���#W2�#M�FԴ;j���V��G�< �@�aL�A'�W��b߾��`��&���C~w�P
m�ǦO�:A�G�1$�O�J9�,k���TYK�%@��̈��2d!3�E,�x�o�-�m|	�%i�C&+k�y�2*�2^GP���F6�"�~[D+C�:��钺i� Җ@�#U�d^���a����
`O ���9�林 ���q��p�<�<w�vw ���(���͡,����G�{~tm�7�2"����F��H��и3z��a��C$-��+�$���"kb>y4�p����U�m�pr޹�/���>R��/���H�����0H�_�sJчu kB���dd��
�b�e�������z$GU�?��ŷ̓nx����_.�d.t������S݈��`���`0	ӽ����-���� ��Q���.��x�k0Z��x?��r�v4�|��ឺ��J���3`J�rx^�o{^C�6��q�=*i�9^�%/��C"���\&��h`<���|0Dk�གྷ�r��K_�}����e̠ttC⎇�>�`�T}[Pi��3�A�X����+��@55�LGO �b��>�x?C]�}u Jso���R�Q��9[� ��,�i��9^a1�y`���5DҸ�.ch�&Y�R�;
�w�2ecf�Ǳ�~��?�a��+�YRRl%��i�e�*W۲=��|�����0�~G`&C���[9�!�	ys������1��F?1�0�xe<�����1�:_�CZ�DE��rY:m	��y������OCB�Ƌ�Qi6�w���$�f5P��YSuʳ	Ɯwi@�#�⺚��/�[�j���P����;�	��׆AKik�8�]��Ax;�x���Ҋy0��L`�W�sQ��H�B�� C�KE(�A��?�,�-�z�����w�qP��	��u�$���4�t��2�/<��gu��h��hx[X�5ʹa�	Nx?�#�鼞�6�Fl�BG �1cT^ҭ��,�����&vN����c�OOO������gum�2� Y�.	���z�
@���C�1
�R*� i�@��vtYz���Kv|�1H�R�NQ0�͸��f.2ІZgoǎa�H�������C%�R1%+���pX�{���<r0�gmb�_�f�feSAG����M����	y(�!�n�c��a��)H�h���˳�,YK�l�`m�c��g��m]�^d<`D��r�O���E紑=zx�QM�x��0dD�Q�UƘ$yxbq����;��E�.A����Q?F,9"D�eCBf�	�;�������*�<�.`�y^��LEl@9� p����pȇ�cϝ�����z��Y7x�1Z�RO���k��5aI��Db����E���%3g<S�屖�{��ݥ�,v�`~�FhF�Ze�t�s����p
�vӤy$< Kt�<�f���?"�#Q��H�e���"�O$|���@L�0��C yMb�g��s���&Q�oW���Y���u���o�i$�'��%��<3i�K���7�����듓�_޼�#c|��x����?Vϻ��΂�l�����t��q�� &�'���1x�x���l�rg����������Χ����9S(a�uz5Z-�򇠻�����_�z������oM�oX�c�peu=<|(�p�M��2>b���+�S�����*��W^�����.��׸U�,�����L7�xK���5	���K)���>=�Mi�m\Y:g�1�.�Ĝ�㣶a���bdo��_����g���.�5�m޴m�>}��k/�g��uD.�L����V���G��Hk��s�e�1�Ƚ\>���96�CE���������	����;��v	�cb�}�j�d|w��C(��Z}�nW�={&?��=lB���|���G�Q[��x���xvo�&��;�h{���?�n��N�>�v�0t���������'O_���imu1�NNf7�Y��:جj;E��[�+��w��]��+vlxL����nF'#`X^_]N�<�@�����w��NN/X]�0�#�z{�L�~�{ӝw�-�KQ�dI�b?s���ڒ�w�}_N�>���W���J�oR��$������;�;]w�MR��&�����M<�[x����/�g�}*�<~\C�3���l�Ok�w�o�����9��ٽ�R��ە���o��Y{o�mN�"��v���}{�۱�������`����0	S��U{4����S���3K#.Ȍ�D\�؉�h(ܗ�ʲb���l��9�b���:�+eCn�UҴ�,/���'O��G����_I�����?�Ο:�E��=����O������T�x���+˫iii����x����si}y-����'��˝L���&�A��1cC���%C�)�zCr��pΊɂ�אoU�0� -�;���8�ݰuٞ�[YZ�n��9�7a�㥱�����^V}�T�R�^�/��OK�Υ��E�l�k��/O���T�o+��ʊ������3u3��!a�s�C�T���%�s��s{XE=�^5!E#|vI�Ƣ�<(5����DJ��6)g��ud [0��R'`
Ξ+�.�<.�0\�+H)P	��0����1d3FІi��ҙ���Q�:��)^q����ϭ&��8g�Eg�`�!ed@����'Q2PՁ��!���#å���$L��U2�4Jț�{ß:�r�Պ��Sy�V�:���'nj;3f�E�dω4�l�Y�dn���E&?`��N"������\�Q�q��v��<��Q�ժ��p��x��0cP���U).�j�M;�8�}x��M�<H��Ca U#d�]Ð�}�t�e)G2`���A�x�2k����oGm8#��o� !Ȯb{�����^^ZW|+OU�62���S��S2�5�d|���\�Q��{�P����#�ۋ��"H���2Pbc�0*}���+*�9Co�'�ե� �B�8��ݿ�Qs���w	�A�Bg`�چ��`�o��Fj�EW�l��M�C�0Ƨ G���"Pr��1C%�����ah���3]=��t�=g5���u�K1�@�y��]�G6�Ѝ��a�F2\�v�U�5����.q*���D��-<��[�Μuӯjx=v�dz����O>�^|�e��11�,�(734x�i ����0��aϐ�7�'�PL{9�yj	�:���,�1�Y�	�9��҇N���3�� ����5��gT�W����Si�a��3����,ίm�^G���Q|jXKe�+j|,2O����4�����:� ���1��T�b��Pex��o��x�!�#w@��%k�e���T}�$uK��=ou	�<�`l��e�|7留/7�)�oN�$C��.i�I&U�m�W^>��NA��/�'�|6���񴸴fm��������Q��I�x5��"�:�U�T�Jxm��#��-,ä��ӌp�D��P!�[�q����;�{M�藪����Sb��o6�v���;�5�9w��S.�G]�h|kkke	iB���c"(�a2>�Ȅ(��Pt�f����76���Q6i�A{LFų|���c�s�MMOe�>r1��x��h:v���iT?tm?���)C�K���fM<��:�_��f{&4������� �3��fI���%y��t�̹t��U;�_Z���y^�,��Q+mn�,V��©c�$y�v)-�)=����d)y�ۭ
���gy��ŧ��~K�����Fm�p0΢:QIm���
teZ�H�:2����G~V�h��D������t@�tŨ�0�h|��N�3��Wt4U7�qC��~ۄ_�B�,�FeL�vq$5$�������%�T�P��dqTF)��H��ʸ�N��?#J�`狀�u��S��L�=|�kzm�����,��O�I�}5=��IO�5\�r�tZ]��Z�ød!�����0"�WH=�PR"�?�!�<c�_A��Ԯ���u��ApS1�)n�E�n�P�|;��v(��k�6�	Xv��T�"�K.��b�O�Mȫӱ���6Ĩ�DV�{�;��-��{�[�����Q�n�� �>�Q��v�$c
bl�@'d��rxL�.Kw�MG�⩶v�Ɐ��P��ۇl�F��׌�k��а��ɢ%���m���������vV�q��Da�(e��@],ңg�H1T��%4�F�c��*J�fdL ���N��G�L08��VG��H����{_�b�엾��}����I�>�lz���3Ͼ���8��W��1I����^WA��(o�2���L���cxg6}����ʪ���A*N8 ������B3:񎧥N����, �{9�/FF��h
�j��|�g�y�C",��1<��1&�]-6����t$�S����6��	�;�e�E�>h;�Cȟ�/��eB4
v4��zf|�cO�ch����'��b`���4��x��φ��	�EU�5Q�i����i��C��kӮ�=iff�3y�-jkA��8�_S��P�W�{�x��'�lqI���45=��&T�f�#i��Q���B
5��8T�u�G�Ey����[o}S�����#���#��5�Ӟ={Ҿ��R||��<�f�Qv�S»Ő效�eg�<���8�����">mK�dƤ	KC�bJ�V]a�8�g���_�d�Cy�w�O��.�s�܍,D	=��ّ3�c����)��e��-t ȸ$lllhTr����7��#4΍�!5��J�\W˰GR �0�����L��c��P9���̰��x��T�y����V¹s����܁�^���Q��a�����Ӯ��yl�: �C����ˋ��ٳ��i����7���w�������~Q6K ��x��.{���J���Mf�K�e�*��6�	rrzƌ�NO}�.��ʂ�&&���K�Ο5C�Y��6(p�����'~#;�)kz���c86bG<��؄�w����`߾CA���� C_�����j�o�G`��$��6��rB` �s{���F��g3-����h
�::y����z]I�v���>+S9�ŋ0k�df�����%+�thF[u8m���gXa��Yb �)B��^�F7߹�d�w2a���X��8S���+i(��䐎���:[̕⩃|����aTm1��Pr �09��M������7��O�Ɠ���䜴�!��yoCH�e�.-��	%m�3�߯���G��U�+c|�E�ۍ��h6?��6�q��c�F@��L���;*�0-Α����V
��a 䥡��a$fS͖���Ŏ��>l����"�X��.��6�"#���]��6:���乆QX{�,nWYG2�ݻ���#��4��+�;'"h�e����ר�|aZO�,vu�����*�FG�#�����v~��܃�@旆c��^}�t1������ۀkj`���0 ���V��X�f��2�-G���d@G0�͈�`E4���a�oKfD�0eV(B�z;�u$F���C/��ڋn�����(g�{1:�6��d�=�ģ��q�hRw����"d�� �c-u�`�&2��1�&�uI�k �9�D�� A���r��?���_��{JF8.s^�u�N�@\�2�m�?xD{%����o"�쾩�64�ŝ@�'�����W,�� tn�lU���Gǰd��gH��@y���q�a���]���0�V ���m'���u���#~1�'��<Ц�xC</)��#	�����@�ϯjc�K��#^۷8�'-��"29�0�/Hg��A����cD`x�;����醎Al�f��
��,��>��S���'��<�\3�S��%;��L�:�Ƃ�p F��j��] ��<����g���ƲrT���%?3-,�Z�#~�=$�6,�dC�����o6�L�yF����i�]1�<f��Ɋ3�4�cU�w2kevͻ��	l<�����Ȭ�0PF$b9�o�%?#��3��9�v��64�Ptt�Q�,ˀ�axc3X5)deE$g{�3���I��1�m�������s��h�џ���?�����R�(���ѣ�x�@�$b5fU������ ��(�Y(���(D�t�]��D~~G:6��D�_|ڶnd$BL�/�;����زE�����Q?�`#~C%�o
�ʲ�2�ƃ�$`��Ob�|���H<>��ϫ۠�lz�)ݔ���s�p�g Zf��v���!�V,��Ay�u�4�g�w�$_]�������D?��F�b[��D#{��uf��][�MhC���Q�u�kܘ�<�Qy���>��ǈDTh7�u�T�uz���7å���>�x"�R��-a@�m]���Ķ*޹�anṡ�1�5�cA�B���y�K�*�r243���aQ�w s�<�gO驍�?�[S� z������F�;{t�؎���E�� H�00D������R�ԛU�H�'"�xn�(R��(0J�E˞�E�y���ƀ�n5rx����+�Ut�C���#Je�#A%�D��𲖊a�����WBP4��B�CÆ�)L���<}/dk\�̠ ��2>���'��$��tD�y:��ɗ�٭��P(�4=��#F36Ƃ4� D]9�<��S�g��F�ol��Y����0x�eh��V�huX��@C��ϼ�Σ�ὁ�;��\���z%�FP�Q'�����OeF��]j���l�K����t�v�̩'���-߷�`ǌ���j�'[��ߔ㹉�h���#<���A�L8ʦX<�y
���5��<� y|��m۵�#A��Ɍ��V
���m�3���E�S:X� 0�"��� ���*�"h?�NZ�fe�����h�s��#7��b��=����^[�>���(`��Lx�o^��Fe�D� 	��h��!�C}�2�ǚ�&��
����:l)H��:!��Nd�*Fo�o�v㫳s����}L׶�ڋ���N�m�_����X��L�55Dޏ�̓��(����3�AD��t��q>��F�G�9HG�(�炒�0! X�[�:*,�(p�q���xv�vfhx�ժV.�b�R��	&�'�C�VCe�׬�.>��rj+i���09�VWΧյ���bxd�9�Y����w��C6lk��8d��itj�����x!7�0*h��s��./u4�g��ʲ�*c*#���#��������&t������ő�L{*�+�+��Iy��R�k4������4��R&�B��|��s4#���� �Uf��Qw"ڍ9�. �[C(��[� r��Y�ńx޶��q�WΙ!����J@�7�ʹw�>{��6�k&+��������R1:QqF����� Xa����:[�}I�f��۔��P��n�j^1��|�m�,�Q��x��꧃j��2	���-4�H��LI�� ����Y��zvM��n�CuP/�6��\�� ��9rQ<}qzf��[z{�2;����1��zu�'۝��n��}R>����6�d����_T�i�����h*ckI�b�%6�n����˦5�"�Ç��W�<xH���Ā���ڕb�K/���q�yqL��䧬ߋ���e��ֻߞ��ֻ�®=&KR��"L5�����3O�g�yFrX��:���'�]Y]M�>��:�D��?�_��n�S���	,�@E�\2�Ϟ��fzⱇ�+��dO�q��]^^�{�<�<�#G�m��fr	d�e�j����"m����t��r��
�>�g�ʑ�ۃ��aY�,�n`e�ƌ��+����<]ȑ�]ҋ��߆�B��la~a�_��=C�����O�~RF�74��dO���!�"�yƓk<2y��Q5|�i=���Ĕ��%ዋ+���kdl����ϥ�{6;��=ų���~w��-w����m�n�{�
do�
�C�2>���7H_�ʗelKJ�cq��k��@�|V�g,�����~��i��k���h�
�PX�!%��|�K�o�'����$py[>-e�f�d�������W��}���?����{ޙF�&�[�P"�1�����gL�_���׿~��(F��ϟOG_~)--/��p�c1�=�yO����:�#ڼ����)cS��c�1�����:}<=���2�Ӿ
�-Eџ����W���E��t|��06~�l5iȚ2{��M�2>td8�ٸF4��Rm9�/��G�Y��
��L�;N���=���?;��� �6#�P�%�ɴ��9	��t�_I_����W��8ހ�V|�!�M�T��.�PˠT�5\�ӫG��z4=��c�O���~:=���:>k�����'=���eY��A��c���1�5͉�'�/� ��h�	�R}/ۣ��w�yGz�]w��Y�#v���O��<%]G�A� ������C=�����ܳ��3-<��W�ϝ=c�/Z|��F�.��=�&c��x��j/k��T<�be�}�����pi�d_]^R�Ey�9��P���yΆ6�5{��cL��J��j=xh�����)D��r�.��_w��fA�H��1���)���~����7��M�gҍ7ޘ�򖷤[n�ņ�]�vK9�g���,Ɛ -腲~�~F8ƶw�o��������3�O=#c{F��S2�^�4Ο{�����T�a=f�{�Ař���./}���ǟLO>������貍kc�?�޾�{��
�Q�f�\@xƈ-��|X��ˎU��3[2��}����h���<}�#���':t�<ƆLQ���I�!���J��x���nR�p�g��7x�t�i���u0Q�#��i���B�uH���䌘涽7g����j�b*���Ww��#<��c��L�ꑇI�+��%X��x+��<����Ӷ�ݔ�l�f���H!��j:{n9�)�_��F�Fڨ�<�<��0Yeȅb<�婍��>�0�뼼����^Q�j;�	��z8}��(���4[��Z(�� ��۾����	֡#��7�hG�8�]�yw�����Y�ff�OR@����4�����-�����k�MW�W�7ʂ�����vxM	�dK"�š`G�t��fQ�f0�D��j�f�~M"�p�,���������������O�'}"=�У�%y�եe{��6`��ԅ �C@���v%�a�sf^�uXĪ`A���ً��&���M��PP�.��R��]>�껇�h&J�;M��Ʒ��?Ȥ�N�~��{W-/ޛ{�F����m�K�v�aN�@��C而>�Ϥ���Ӄ?da	����D�e ���'i٨@M:���7����2�����M�|/��R��<��)�~��?w[�@q �;�Wr����~�0������fF6d�7�,*3ԓ��^z�e�D]�ǎ3��`\ �а������0�0H��@)o/�\F�bx&{҆#�ʃ I'��Cq�x<��~C� ���m���1pv�2��<tuD�����-t�;�U�fx|ꟻ<�Nl|�������Y�J�z��IylMH��ųVI����T�yn �����nȱPn!w[&B&��� ��Q굾�5��_K2C3��!�gTI���J�"���w���4!�@5<t-��zU�3��� �" G��xcQ��943@z-�F��>Ȭ
���M����'A���UŅ�'�oru��-���MIY��}~ą�E�0��B�B%��,��m�uڱ!�odE0��,�}���Vh30J�*KS3ӽ-]��x���'x�_7 �Mu���C�2��>>� ]��f���D^�Qdב��}2��`�7�%^،�P(:��cO=���+����x*���5d(��'�4��n�N���Um���ĉ�&Xh���"Yz`
M�����` ~g�u!�1r�͢�hI� P��(KpaȠ=�n����糸leT6�?S3�i[�c���6ۨ*�1O(I���^��A3���ch���vYlT�f�I�x\ޚ����������H@L�+�F�؞>y�B�L~�w7,{[xE��s���8E�'^�t�-(�D��!a(K�v[�p����ܨ������w�!hx�n��|OIyK�f$\vIp�xG׹7�{�v)�ޯ�����&5�1"�W����̮�߅7-�eD���)�˔k�MM8�W�Ӻ���$#_�Lk���5�������ݨYB�C,..�^�6xbn#�W[�(� 3h� ��aɌ��"1"��o����;�3��Eϝ_��j�ˈ��&�y��Y���21�j�h����x~�l:�`/��C�
��� j��G�p��xD<��UX��n^�@�|[v��cs+��M�x�d�喟pl��&[��6 %�ml�~hc���f�-T��j1�7%t��4�@~+��=GC^��4����'N����4>:�}&����:�b���l!vaa!>|؎���y���~R����z�['�����S�Ed0(c�<O���}�E[���d���O�[�����~���_�BZ:�����)׈e������b�G���>&��'�z!��Gf�\����^=s*��o�fz��MA�n�bV�N{�7�;�+]{�w���Ptl2�3r� ϼz�^:y�����[6` ?�P�L���f���#_�q(��"7m�!Xh��i3�Xa4�}SSӵ�ɉ�޻���Gy�g��1�))���Z��[���[�}�1E����PB�G���S.�@�����у&&x�LC�z�Gc@��!�LC��P2�L�܈��0��iD�����c�O�8Ƴh�x�چs�����@�zϞ3�_�*B�Ȣ�Ч�Dì���/�W�x>�e��3�~���_��6ʠ���tb�p#��dw���1��}&�^�Ͼx���ЌV6q��m��-�ބ/No��6�Hh�L&}GR�: ~�3��h}|b�Ӈ\����_4"C�0�7]�o~`s���N�}�*�2`�Wx1�gaFX�@�&��1��!H�kht����
��`XT�T���@?Bm)Ȍ�@ �B`����� �8`�U�-#�΋+4.e��x���8�vK��0xd�kb��x���ƈ�ؤ�ڬ�Q�rtf��Z^&����(2�<y��q�9�!�{�λ�)Ϛ,�q��V_�&�KY.��z&ӁBcll�w�9r�
�X�!�_�E@�O˫|�^�~J�߭Jꕡ'�`��OƼ��t�W�!��`|Dç	S�LM�����hl!��&;�Pԃmc(�$(��7 f����O�.� �f�H��YQԅ����ɤqn��
"/@�e�6`�%S&���S�2lq2O��8�7]&!�����[t�T:�ڒ]#����2Vu2�G@�~[>%�������P�Ȯ���7�� Q�d�����U��?�0���e�Co,p)^���,�"EL����:C���b8o��-��
4�Kcz�tN0~44`T�QI���$��F1�ztF�1�=C�~�s�k���B� �_ĥ ��wl�0�A���oW(�#���N���l�Z#G�͎�Ηr�W<^ ���@+腱`N�҉�:�yM�ۃ��Jz�>ґ��@6,����T���¯ɡR)�ȫ`� w�a�O`��.Cy ���(���"h��Ęf��(BG)�5�#Õ���of&,�5!��cuPw�_�CG� m(P�"���j��G��=�M]2Z������?!!�����x���,�H�
��1p � fP*ƍ�����QJ���QG���z�ǓifnF;x�|ɇ11+4�S9&�x�0{&&�)���= ��)o+*�t�,ޏON��:m���@
����P�@����Ԃzh[�%��!0�� ^$��Z�q��L�1�1<ҸrNl���\z���1��)��tĶ-���U��G��/�\h�L�z=<`���"�6၆W{��a|��諌�+/HG�ˣk5�7�@�<����c��4����@�����h;�uB����'cdb������%=r���X���t Ɂ��xFd�%�1gdHت�@�4�)ʓ�YxH����E�0��,H,x���Q�5
e���VA�9�RɈ�5C�a"�IN��))�QPG(����0i��!!a��J�)�z�֏�Q��gó���S��~Ǿ2C�x+0��<���c�"�Y�z���S�E���$� � �@�=%B/�̣2q**�H�0�<��x�h8���$/�}�eS[�R��pk�_��.��,/[�-�t
���%%���V*8��-̲}E>vg�:4��@�ײ{�	���Kn:G�ރ�611�B�A!<Ι 0��|��ߐ���\A�:< i� HG��Ȇf ��^�<`���h������ybxI� �;�^�T0��"/i1&�2~�t<�F~�\E������ǆ2`�m�H������D�*j�\チ���:2�a:.�z@�WU���)B�R���(����Q�U��.�!�/�K��N�A��e��vgJ���z��B��#lC�j2�z7=�gZ���k��`Ix|�
d��xh�7ҕ�o�?�[��d�|_lbl4M�|&F�R2���B� 踏�k�#�fԼ��/h��DN�B)�3ɺnϼJ��s-�~�B=��M��7��2E�K�A�Lů�u��h3�A��.(��VE��I�O_�	�r�^$3��;������3�����Gx��<�\�,l�1��w�1�!A�/j��;�]~Qܥ�t������m�"gZZCq\��4�����W�F{�C� �7���dÕ��Wx9�H���du�1n�Q�����2^�:"f3�e06)�(�-���0z���1�$�٧m����0��dб3��4����l�,q�	_��iFxy��9+#� l�e�ɚխ����è�*bG��C�y�6Rp�sB o��pJy���<�{�OE֮���f����Wg����=e�C�s���J����
�)A�eG�YA�&E�z���!�t�g�5� �����1T���S��U�ʭU4�Fz�)φ���-�.È�C1���Ĥ��@1��2&&&��^�'qK@=��ש�x(\5��dO�wR~œ
������3�e0(��&�y]��е��b�"���a3�</�������^1�:��� �)�'���GՒ��}Х͎����WW��7C�U@h��S��0h��=�w�I��^����%A�V ��F���%��L��x�&_�A@B>Ӵ��l���K��F�j���X�#���]��⸅�=��_�#�R�˫GK���~)O��!�h	C�@�e^Sr��+��?x8�ݿO�^4DWYz���r��.�M{0�� 0,m�،�R�xb����l���i~�n��`l�������K���x6�^@y�|s�PD���\:x��γ}��ċ\�y�L��D<w��6�G���0Y��l���s<��1�?�kC����	��Zc�\)�������h�j����14[�V?Z�m��ιá!��@���"a������	��9����`Ua�EH��Fz�]1�q5i�ظ.��K�[ޜ�g�L��BH�PYy>K��3Ϥ���jZ<N���I�E�m�<�V��lm�'�n��N{���R��3z:S�3"�E���3O>�Xz� .@ѿ�gҦ:�$����� 6N�,���Lzǻޝny�>��K2(1{{E[r���+�_�|z��G��ںm�Bv�>16f� k���tcz�{ߟn��Q�L]�3ؗ�$G��x���ӧ�q�Eu<��|��o|�ɄiA�d�6�S������`�.9�` dI��-�)C�|Ϗ��������/��X%C��Ʒ���V���8���f|<ը���s���'O�Fm�&4Ζ�^3BP�<3 	������W���ѱ	�;Ҽ�q�V�3:��R���H��}_K������	� y���\���{���}�xz�?��g����T}����������/�o>�@Z_Y��0��W����ciueM�iW��� ���԰,�5f�~��یҹߊA.--�����J_��ӹ3gM���%Ϥ�s�6���O~��o}�չ���cTʷM�xe�#�,�ҋ/<�}��t��I�(0A����_��~4O�7<�׊�a�a�ey�i���yA���O������NNL��{�L���1>���$� k[��(�#=��������=��x�!����������m�����.�U�|f��ɪ�~3��9z������c/�x4�z�d:u�x:y�X:w���{:�=`h�X�@a�8]�p��S�/c���2[ǬY��o�*�<��<�v(�4�.�D�1��6m'?n�1L��F6�z�8���O:���)3oEyx��aT���) �^�PO�"T�TH�!/�����{��<�f��+��rN�=�r��������0Lf�
:s#�cyâ*���2�X��G�)�#a&�a��&�rЪɳR�k@G@�n����T�`RC �P�ьkb��;A�������4�#��	�f�A��9�G��-`՚+\Y�7,)v�]�ɪ�m6ÔZ <���N;� �s
2`tt��ŀ[t�D<G]�`o��[t����nב������'��ɝ�L��	 9�<�P26�⋉iy(tJP�ˀ!-�[hK,�0����û�^��@�mk�0�4�$��O��0 ��B�3����P��5���7[\t�C���C�&��v���� +���M�0���3�za�/=�3�WQT�7Ҋ�{��F��y*om�� �Q�I'�Bş�L���⟙)3Td�z�T_�\\���...�S/�?Ǒ�e|
oD��#��%λ�O���M�)�P���m�NY�gR��pD�F^�Y��1#A?��X�n<d&㛺��g5�,^��qC��Ø�*Ë�{�vֻ#� F��7f���7+r���{�D��	��M���if��N��-������Ef���K�4SEN�^���!^m�Y�����U?��;F��1�rɰG(�k-L9�:�X��l˩��KG.(T8��=@�S}��C�����!K�F�O/�� �Q7�`�Icv�wC���­9��ֹ-�(�r����G��N���-2g	���N8��"���^n^��	9A��<��f�,���[�x&�v����Qn�s���x�B+�F�u��_o���}����p��tN�O��P�A��(.����,�����xxhlt*M����־�$o:/�G5�.��r�f|f4H�zQ�%�(����?�_K�k�iM�����D�_f����9��Æ�dX[��ވ"onw%�������ɨ?����!�KQ������aK���˃b�����8t�[�0� �Z���nK=A S��f����G������<Z�k($v14����Q����X]�.p�!�M�,�x���AL���N���i�.��[{۵˟!?ʩ[��� �ę)R�ꊋ��L�mcx��q���}���,�G����
a�Ҟ���=�D�[ޚ�ʰ�k���5y	�`UY����Gd�u�ѓ�h��gwpXȖ5��]�S|��Lo�m�2}���ЙǕ��q߾�O_��ZY�)� �P�2H�	R����1$b���E��W���zy��4ȓ���b����z�"P��75$I�<�651���S�$�ci� 0p�1Āh����6��q�����"�Y���;\�شj���[�-?�:bƿ���n<��4v��H�&Zd��#��d	�ظ�¶|щ�QY&aT2T��
2!?�x�F�&�ڨJz�!@hM@�];������:P�m��-.�!a(�W*���_u��ְ��Qo�+`1 {(Z9A�3D���Q�Ex��̴�Ҭpr&����;Jxw����Æ�Q 87@W*�ak�i�����c˾�R����'�N�|��FՂ}��o �Rq&
i�WJ�J��[�M�^<�X�����(�A�(yP��2�0�'�g�7�GC�3��Ec��Y��)ތ����*�[t0Pbh��<5y���k�9�Fw�"�͆���ɒmf]�k���^��+�s�F���Nuzٴu>���!/��2۾8�a���{�7�Q��۹���m�h���x�	K�
i0~�+�")<BB���Bz�]�9Z��8������.�g�Q�[/0S�0����^~��t��R kf�by v2#@��CG���o`�T<��5o��#k]O<�p:�ҋ��_�iwN$u:��o|���7�9�x�-��,��o��£0{&�W�6c�������/���C�'!?�d8��S����}(]����,L�2�p �{���ԉ���C����=j��rK2�<wf@f���I1��-�Pw��T�����O���u����{��ޅ�.ھ(9e|���{67k���4�@(,?��?n�[���P�:�Ćkd�e�͢x%C.��D�eC�[��7Rr�A1[c��p�����,N:��@b.�,	xH{��=�Xpzjք�Q2��@���͗���-//���=i���cU)�'��eLh�1%���r��1S�]����B-��C^Ή�8'/�I���-fU�M~B<9�+�nv-���1k�,�[gґƓ�B��5l�y�h�GQ�>��V$�ٛ�����F���>��k��ٻ�Я��5�I1!���Ey�ۍQy�]	���}U72�S�1�3��#���L0�Ȱ@9�.��1aI�P������a��2�׃��G�P(#�:Ʈ]���(�oz�긥���y+�@���g��w��C�x�Y��~Q��=�L>r-�Yxu ��uv�@�� �r�6�Gk7�C�'D��@G��^�W"5?N@^гgH�Y�)�0�T�8S���3s�?#χ�]�z��tq@E���R\,����Ŭg�01��F��#	Xj�=u�{H8ڛ����5�n^�oG�@Ң<DG�PPjO���x+��*^���X�`8G���'kC��/؇h'q�ؘ���7��S��	ĄŬ�ɀ��Ex������aA�d(㈂�!��S:2d�7<'G�����\B.��9S�ʪ�& r@'ǩZ���0d��Ѝ���J/�H���'߈���1>1����׭�Iug�ٚ��b"J �v�dȹ�� H\�;�u�=]�t��@�p�i����N�@�=��`LF�N!u�u�W����{t$�r��(Hg6l;��w4\��h_3�@�2>3�^fv.;�E���=����*Ox�Z� ms�T�*���0,����"#�
�F�g�lybм�t`�pt$��|�:���k�2ш�T!�x{̕ټ��s���y���>�ӉE��F:�lbt��[�0��)�.��޶қ�kp�^e�����y�L� � 
eM*��,I����Κ�o����#hKBf� Gfq쌡i���10h�n�/L��Gd&i"gx7�?�D{�a)�g�9d�x?<���G��O��t̃fm��kJ��F�c4A���_���KyЮïh�Z�����fKn��|�\T�ȵU��D�M�@[�6.\N��Xǵ�����/�!����ab�<o��!/��$0��a�D��=Zh�(?�>u0� �(�À54@�ms�D�m,{�5�+}�!���z8�1h�hF�?b��w%���w�h��B��#&����up,;���0��e���q�vTG�?�J�5�c�r�y��>D��(2�����ٌ�VT^\����w%�f�o�\�s��H�e����MM��Ta�iq vM���?n}�#�_4-&�B���P�!6@(�<.4�Y�9�
F�Y[EW~�`�<ই�FE���q��m��+�-Oԥsx���7�A�E� �۳���>��p=��s�y��Z��?_��͗Ц�a��|���>�T5�ݘ����&(��7 ��%h�V��K93d�����m0ʉ��� �$s��7�����9X����O�Ƃa���-I@0�@��@YbזV��VcFu����s��Y�f��h�`�w��
�u$�3�^<�F\A9v�������B��O���J���iK�~���2rYM9��]�q��^m��YҘ �S~vR��r�,C)�ZlWR���=�at6�R����g���TO�8'��.�Vϰ��c�x�"�I�w��}� �Z����[�;ȏvif\aé:Z<C��uɗ����=P�c��2_&%6� ���4H�j�ݭV���w�2M��&���0���1��������IeD~�
pA��#Hf� C�E^�"P�:�V�r�,���� 
Fev���Q	���a0^,���@�ÌP�W6f��H�����uދ�h��!��`�c-��A��8��=��c���j�������_��"��td°/\����eޟ��]&y�-�Gh�ՙ)�����0�S�Q��Tu��&]��j��ё�ߚ�����ƃ'CA&�K��!�[�_�D�<k8�[��=gdL�WM�%�U��w�3Ji�V��:^ʶ@I0�`����9'"p�����O�ؓX�Z�RԐ��j�'fI��ݢ����hMhuJA!`D'C��>�,%�)w�����4+e�*�W�0�����g����#^	����`�d�M�@�R�{�<�-���6*I�|��l;���X&�7����F�h~�>���̢A�S0umFB��*�Zzn����X��,�7��rn������T[[N�چo,e6_h���|
���t��A�=BIL� ?Ñǁyc L���b��0˳<;���Ϊ��`�����h��cu݆:�pB��g=��)d�ԣJ��y�%��W�ޤ�x�=u�)۪���j��ic�\�\]RS�n����4Cb�0�L����y}�	��o�^�[�j�#�d�2�}�cG����_�49��]�� ��c�� E�uΑ;Ft0[�U�f�eI�ޛ'$�Oa�X�c�%����.�K���ɭ�]��S2�w귂�:�p)������U�{/[���vu�;dD�ieձ1A
0��~�d����8d�����4Gi��ި��~��S�1z%���A�Z��S��溴��[)>ąa�h��:G���Ey<r��	�&#x+5P�鄶�@Ƚ��tk����e(�'^��Ŷu�B6�^{����s�=g�E<K/�=9'Tx�-��;��^� h�e�-^�������a{y&�W�953t���u�A�q@�r��|�_=c������y;�Lt{��u���c�������D#
�2>	��ju���C
-�tK��n�ѓ�}�������	�G�Yh$�j\,���6��8HQJc�`����=�;ߚ��X����f�B�3Ďi諭���y8=��#V7÷Ŝ2��c늊�� ��oW��ƛ�l����9G������}���?=��#��5"��h����(�����g�����~_���|�I���[�ˡ0{fB$*R;���/���{���mxų��#���i�'>���g��M7�t�Y>[�PݰM�^�#x��'��=�N��ëw&&}�%J~҉�ˌ�]ጿ����~;_��C7|�/F�_��ܙa�̤����c�SS?93���W���k��{j���7�{��j�^�-��i(bx�\�H'OO/���y?bG�+�nt�`[��1� X�[p7�Б��?���{����I:�˖�e)PIS�%3���_�ڽ���@ ���]e�|l��[���J��G��w�m�Ψ��I�N �s���U�n���?����7�~�{Uu��h�/���wh�;tM�c�ӛo�KJ�Ұ�0��ty%<[3n>��O����>���M�N��z�|�cBC������O���W�J���[3���3P�@:2�8���=��7ӗ���t��q�i}�T�leA�y.Y�����2�'Lt�[� ''����]w}���N2<�d}�����������ss�O|�n�!��a�P�`��Ĭ���=C�Bm�e�eT2���\*V���Elё7�G���b^{�CQ��uq3`z�0$��8J	2��-�4�lSq�����+"ڊ]��A/����' h���Bx��e���b#&O��R}X.mw/���L�ԧ���N�g�w�J�Ksx&i�A<�N�k��^$����Xax�m�ZGF��SgĠ�ȧ�-ɕs^�n�����i�����|�U�L�چ��'Q@U˷΅�P�'^_vvfy��0�b��?0� T���� K����-����#$�#��ϻ�XZnx�����+��Ф�/cC�@��-�g��'ߩ YQ��8���A2�2�`Px�fmC�4�F(��t>���n��;�P���Sb$$��#��TF�[�(�'
�>q�dA�����Wx��kd�p�����f90�R;E�Ϛ��M��{�Ӿ}��#�Ӯ��4�^33���9��+��d��t��k �<�K,[�����|Ϙ���]2��:0#����:#�,��ES����[:�76�j"��(��:���:J%b��a(�k��n�]��Xϲ	�BC�=�/e�DC@,�3�|(
�"�����
M1��l[��*Cb��b���pP��㜅]��n�bP�=q%Za�<s�?v���C�=�Bqᕀ8'(篝+�2�v���1������)/���=β���&_������af缴h��ٴo�B:,/x�ྴ�.��M���M{�g҄� �1�X��ꉺ�.zrS>[Ȗo(�� ]z>���9Q�d��$�ͨ$����+G̨㦁H�6�l��]�9�b�h�'��hXU�f�?����(f�� ᨈ�>p��� y,�l7$![�7V׭�R@�g�*�#� F���q��Y����>.�,!����l�lt3�G�.�L�Q�%%bgK9����Y�,���4���ӕ��`�DKհ�b��S�ϙ�s�KՑ�6��޽�Ӿ={���kN�v隼�:-H<���y7H�t('�-���m2�Ei���amϼp���2ػ�u��ё���б6$ۈuy���={V��]b؅��Mf�^�8Ǜ��yopٶ%�&�2f�$���DA�2 )��"|ц}b�O䦶�-7��/��=�S���۳R�MP�H�n�341Kc��B��,����`��߆{��}*˰i��2܉wJ��(0�o��ç�x���2����[��9)�����Iu�
7ID�prΈa|+�-*	B��f��#�@����#�C3�C�Ȉ��}Y�w�R�+�4Cy���CH���>���.�0�0�N�_�i�j�fa�0<�E\D�8TO0�C��j�x���� o�����#�Ä����sBU��k�S�THؕ���-\4����vHBv���i)gܔ/�J5ʯ����2>�6�l�573J� m��:�`|n4�S|���*K�9����i[���vdD|�K�v.�Z,h�a�T�lTZ���	�;�C�	c���`Y-�����z^��Ďx'|1��n�����(A��;���B�>�Oн5_FgT�� 9����/�y��2U�:��&_Y�qc�����?)v4> ;7� �z��8�x��n�%Q�X`�c�?Ʌ��@�+m;�u�Q��Ɗ�W�v ��A�&P����xS��o��lߚ.8�B�q�"�ҩCyX��0:Fߍ��5�4t�nxU�bΰm�K�Ykt�FUʐǥ^�P�{u�.��ʍxd<�ա4:B�c#��]y�8O�ׂo����G#:'V���3KVx8��:�[m���P��F�<-g�E����9��?�s�#@.�'xu��Bv4>Eb�l(�	��߁������`Q=���Q�+���[^o1�a��n�
_잜I�s���C��|�F8�:�Ɠ�S�(A�\v/����Y�D
��� x=���<�({�ԫY�y_�F�<�2ì���Y��Y+^�]���*Fx0j�a7��c6\��CAx�*df��tS��gg�D!o�a�D�<����t�ф��P:�A��^��,���,�1KĦX�u{={q��zA:+��[G�����Uޠ���n!d���{Ei�|�����p�̙�����67k�լ�UI��^*�(kF̄x��ٳ�ZO��-�CO��G�Ll�AXUy<(e�q��b߾}f�>T"`����Xs�qF���^�Ⱥ2�%�)��N����r�7�tK:|͵��. !� C:1f}s#=������3v��"jʑh�bS��Mx>:x�]oK���1}	���3��z�����S'ғO<�^y�%{�݌&ڨ|ȋN��]����nK�v@���h1B0d�V>�*���/ٗ07�Wm�4�mF�ő��D�ګ� �%���]�w�1�c���M�\·���佚$������������?~�P�|�^o��b�;���a��/�X���*.	F���<`T̢t(��6\�@^��D_<(Ō�[Q��(~���x;��a�iϔHQxi��(My�ا+��f?�om{�Q���Fh �j���>���&)�}���A��a�%{�BgE~��B���&R<��!;��m���	x��G�e��� �!mC���GFˎY��!G�9��r������<n������={v���م���!�)]���������Q��x�ռ	Θ�V�0��L�9�22,�%�"��8hpFӖ�4Ι�l�0@�a�K\D��,a�A(�F�k3�(�f�rGt�<��o��%�6��>�9��3�ʆi�I}��C!�6`r4��hGD�Ν�6d,�d�����h��������z�`�u���no���AThuS_ԡ�l� mue����������p���"�J�ƚ4��@��4K�`CH�g�\k�ê ��2\��/)���*� ��'��'�w����=�a3'H�,�y�V��������.����Kb3�)h��ȉV(�#�6��ɛ����kۆW�%�S�Pz(�R��W$.�T�����,A؄IHl�э�@��I6�3����'>4�5�g����A��"�*:#v��<2���W><���	K�VU�J4�z]���G�Ñ�ȶ�!�t��;�Y.�t�(/�b��Ǉ�u�a��+),�d�-Ͳ�7M�1x%3 ��v�ߚy>���d b��Z�s�芤s�q��"���,��@��0t�ǌ��<|Όóa\ixSh�x��$%[Cn&G�������e��+�[�CX�,r�,/<���]��	C���9��-0S����$Rt��*����z)����v5΂��������O��1�.(�G���d�
n ,]0������R�=�.H���I1��VU�����e
�Ak&��``���0�� e�}�.�[ẻʸ�G#���g�<�̙e�A�:��m��ձ����H�I��p5ޑ0n�4��E���*p�p)H�|��`O�E��<y�B[��vH�a}��N�R̆�^�� �'�p1!�!��^~�S�ǌC��lb�T�@9�V�R���:ڠ��g^p�8h��T1��a�V�9��|Z@^~e����~�R�`>��5�y|��k ud�:�J��ˁ�O�ZȊ��s�x�8U7��֋
�,����,K\����lH�Kb0�N3��(5h��2���S{h -̣�l�a�A�X��3B�6S U7B�GP����FA�����A���a��$v�<f`L���\�� V�lg�`x0��Hfh��n�v2�����s��܏���2��U,*��.�1>��S��m�j�	jkC���O�G�<F�ق^k�9`����$Pi;��֏^}���3F>ʌ*:z�X2����=ێlڱDZ�+d�o�V�^�6����6*��62�ቂ~��K�m'�fm��,��B�@g!-����k"o7�|Q�2`G�J
�įFReG�:�� �����B0�B'���ޙ��|bFKݩ���P݀Ŕ�dk~9�K�`Ɪ���A�<�\����5�!Z���=��8\N��������o[�����h�y_)��&�L��5j����ځ��n�ϭ�MK���+�z!�a��R�:�/%�� �{�eh��<���~QC���ml޳\�����=XDS�ީ���� #����2�os�θ�H�#r	� q� `-�w���!�o\�d͍��"�0�a1`�7m���� \,�;4/������p�\.�o���Ծ2�0CY�+����<��u�O�M�U!��;R�a<aH�y#4��#��?B������MM�kfoL�NlUY�LC�`�_�ߩ��b�Q�w�0D�7-�+2��P�an������y�.�G������҅�� �V�Zy�o�7�_�����ߺ��A�Q?i��N��u�~zՌ�[&@�w^���ˁ�A[p�� ����Pv���G��8,��oD@M��e`(�'3�tr�����jA(5x�Cް���b�B�q1��q��4���6�!=_��������P�v
���7���N����=�g;:Ô�}�<��y*��B(}������Aw�y������ ���$���]	�
��P�Ɣ������0��uF��
�U�������+�X}�c��٠FF5��냘�3^)ZW���9�Ы:�5�����aDyC˟�F�8���� ����}�
�~�_�G��� ۔�t1��0�8�� �y�b]-��H���jS�Z��ԥh�\��n�uB/�;���n���y�n�6
Zy��!�B�4���F�(s)�_/lGk0m��a��5��5z8��#�������c`Wx���]�����Np9<��[�;�#�n��`ؘM�\k^�q�?n��"��j�������Z�_�&@ސ��`z�á�A%ŭ��n0�v4/��y��z|-0T)Ef�B��l�D���Ac�H䋲�j������?�m����l!c|�v�3��+2���$�&�@��ow%�/y�9�#f����C�"�h���U��\�0�BY�v��[��<�F�s`��ö��0�񭮖˭n{�����zBGH<P����P0��@�G�� ���w��7�������h��nҳ#�Y��R��8�|z��K]�zvBx��?l�|[��$��K ك-2on����h|"\*v�S�b��W@@(h;C�lG#��L�w����h\
�ϑ߁���e��c@�|���9`��� �]���-����!���)@���Tf7�c���� �l�F�A��|����u��sB��(�z��Ȑ߼�b0-��E�a��_y�/Ն���	.V>W/�O���+���jE�7T�Fq�O���R��J�c\��2y��H�ϛ���A��iq���� y=��N�ڮ��0O���G� ��1��E�h{��Z��}/��|���oѨ<��.��|:���v0�u��#?��@��5�Q>u� ��by�V����<l�������7,\�L��M6��=�����|#!��۝�eE\�ȵhh��ky!q�"=`��0<���ȟ/<�y@�< ��������H��y��q>xzkϥ :"4�	��^x�{sjj���*�|C�˸��:�;��6x��y��a�|��O�������#};����<}�ߡx0ҁ��A�.=��f |]�y9���i۝G��� q���o^y�*��w�k��u��Z��>䙺�ǹm�ʥ4#�Ŋ|'"��h8�Q6/ ��&Ho�wځ�o�� ���<���w'̗��`�|Z�/��n���B�����&uK³�q����h4��b�d�TZ�O��b������h_u�#LJ��̐�VB�*�9�u�A�F�՞z��_�����*v�E |G�����3�^���|#�{�c�|T�W>�:I�Cz����m�bY4�A�F��*|aF@���ʝ��0�aбM�Nh�;�F9�x�'��B�/U���1{Ӫ�j�P�`|���A�މ��Tt��>�����ħI�"(���C��j��ʍZ�fD�[��ym0&�^ɻ���{�M���m�!�˙�B�ccc�3�����.;߮]�D�p���|S���F4�?P7���;�8�M j)�I�Rfff��sZ eaA��$���'�� y�3==mG��#e��z8�v�>�E��	z��!_���%~s���D:m��}h�s{�l�oe�l� aL�?����z����}�F��\������Ȅk�C>��C蠿EY��s� ��N"�I>��&N
��R�k6�;�*jv:�c�b�W˥�oJ �TڋbW�&&�B��0��@���(.�e������I�6brj��O��{�(5�r�P� ���DI�S�lG�b8y儡�QB��h_����vV�(��)�����՝���r�[^*j�т���~1�0���u�·�FG�o<^xBdD>x��q�s�h��-�\'��p��	�?���I ��9�Q�a���H �v�1�[�S���X�������bnZ�t>)�8����x"��L�(��1~���imm�+�s�޽ی�O�^uC�9��єŻ�����7ub�"t0h���4^�M�0>�-�xK-�ǧOc������}����m��'�N����+���!�W�6L�|7xaa�Ҡ���n�a��<!c��rYZ����O�aX�M���e	���9b��9p�έ��u��6M�tt�/�yx�R�{�����e����B����kkccbl�XlM�ۥ�b�=�n'���H^���~5F��]��9��Q�0H^.n����^JO^YYI�����}��g
�������w��izf҄�oK��eg��A:��P�Xߣ�>j����wR�������t��)�?7�+�r�-�w��=�hR���3��2��ڦ�{��_�|��ߝ8��R8�!±�_I'N�H�3S�;�iff:ի>lNHqO=�Tz��e�c��7��8��>}:=�����0���5�\cFz�ܹt�������{��/s�u����Zz��gӱcG����ő<O<�D�H�Ї�M|�~�mo��NH���	p<~�x��7�O�?�|ڻo���{ia���x�7|jtt�e��C�e�nTI�Pػ�F���h�<���cc����_�՚����_�����O?+#�E��-�u��%��4y9&����a m~~ޮ�$z�����&�a�/����vJ=S�}�oS=�����c�=f�Jܳg�!�� �~�����������MigΜ1z1FMY����q<���_�����,Ґq�V_����g>�t��Qk����6�c�u�s�Τ�_~1=����|���瞳����_�����+�?�������,0 /O�#�.--Yyx^]]��ǎ�b��'�;�&/�Q<�1)������/ӿ���>��ϧ�~�/ZV��S�����jx�ey��Ɉ\���gB�rA��F�~Rv�A1}�H�RF�!H�����w��]��;�bC �GoDp�k��k��葤34��/~����������[C�1]��_�%�5�]��ğ����7�`H�?�h����m���r��)ş<yR|��C?�CiA�����'��:g�����|�?�n{�[����G�$厅k�+Rރ鼔�*Z�?����F����#��G�#S�x�S�OX����;�u�x��4?��d�����������\>�6D"��A�>�>����OZ[O�>���qq0^�2l�F�Tdq�ϲ��=��#ֆ�����tm9��[o��|�{~S�6L	������T�76�ݟ��O�k�Y�M� Bfya��G 2���b�YX�e����Ȼ�?�A�歪j����{���v�n��F�����^���?}���������������������C�>l���Ï�p�K�����Q�N�K/���v�W��ߞ>���7�'��r��6M�dl����n#���_Ҍ��n��F���W����6/`(�K����l��Ǿ?���[4:L��������ҿ�k�f#�G?�Q�ƴ�t�{�ɧ�o��o��}�'�����Y��}����O�|z��G���7r��r`�K{�����T���3طo��7�閿����o���^b	���O}�S�?��~���#��}���x򉩇yd����i|b2�ٻWJ�G�ߺž��RA��Wk�.�{��4�ayJ��hRp�}�j��I�\{MڽgA��wf�iM{������%�Q�)���>��o������c�J��:t�<��ӯ��&	�D���+���=�kJ�}"=��#����,�o��o�����M_���d������B���|�y�4#���1�5�?�����cR,A���41>e��_4�O�xR�D�]_��cF���?��k��C4pL41���Ld�	�_���g�̟Q���l��O�^z��oZ=^ߢ.qbC7*]P/����u)���Hem����]wݍ���O��e#�5>@���/��/����������ߚ������O<i1�]w�e=����g���reeم������4gμ*ݫa�F������S2�������˔���?`�
#"�qZ3���o�Ǜ�4�\&�幈��ў={M9ē(�Voh��d���6.��.�i�![J{���ԙ��z|�������������O?��������@#������l�v���
�	@ba�2{ՑWU� #�y�M�ذ���?��J�/����[Yd�'��O��+%�6����}�2���x�-O�㻬	Ǖ 5�,E��
�R)>�Sx�Č#@��(�9�t`$7�|�	���z���&�X��G#�'N��M�5f��*B�9��V/��w(��	^����H���B���7�P��x��>��c�U�Գ��C����/ڰϝ�'�zF�13l����y�3~�-u��KG@.x@�/�	�C����/ir�YOo������ߓ��t�=�o�ūf@,� ���Cx���#�#��hM��GL��ô��j�!�h�������ޖ!��e5l���P>���(���?�G�H����!���|�G��0����0� �C�,���I�J�>4(�"0nz4q�1@L܅�^����x 1	�cp������B�;�ӆ�7���6i��Q����t˛�dF���Fh�!E��`�����M�M+�$���m���2$�ŀ�E9�E������\#/א�K{0h�W�]���=��5gxÍOB�c2%5�^�F/�w�-4�a2z:
��"0�!�ݻ_�B�)�)G�54r/xiqń�h#h�A���R��qw��믳��G^�_��P����0�!�9=�+�..�f��*�,��Q����11@��g5��x����s?���������_�o����x?��b.�#��f����	;2��0���/9�����^�'CZ���VW�ӣ�<�^y�X:���&<������bX�2w2��N�x.���PO��"7Jn6�I�񽮰�7>@�#�Ez5�A#�i�.����0>�������6�ɛ�@�O�'k]_��WL�Љ�:H�>OB@N9���c(��P(>�<�,D`X�^(�#F_x4�$���^MJP"�ߕ�5�^����� �����t)o��ƨ+"f� s@������3�����L�$�\���8F'����0 �9���1��2�ryD)���OB,H���Ɓ@J �c��4z?�fa�`Hv�7�!`b���9�co6E>�܋����,BW}�I�F��cx(���x�xP|�0�0b�(�7�����gM�:GCJ������\WL%��h�SO>��ƃ�B�M�_^Q�H��Η^y��1������U�9G���Zq;R����%�����^�6��o�F�]���Ķt�������i+���� �(1|�� ����^Z^V���5f��Pq�?�����ȓ|D�B(L*~�G~$����׬��/���;��;f(������w�"'�Y6 A	1���eS��{�,��pO m�=]f��=tO�<n^������X��;��zxJ�CEMO��%w3P.�Ȉ%�/z��A��>�)�m(���M�@��1��a�ajz"ط_�r��N�~��gu�n�Ҟk��VuL�xF�ː�0?�P�/��l[֠��?���?���`ޙ�����6l�7��(���f���~�����ȑO}����/4⼦M�n|�������~QF���Fm"���M?�?a^���ݿ�����&8�1��\�w�,���13̡(b9z9���%���+�l `������,e��5A?��`�Fy&HĜ�N�k�@��N�Ar����̑��̌1^��9}�[����1:�`�N9��OLh���m�Cΰ�L��Gg`��7#������������~��~�:+e�2�R�Ɗ�`q`GQ��?���d|���?���]�;�e�lxÍ�3��������������4�"ʏ�؏���ɟ4��ʯ���X�����#$C�5x>&���KV������J6Lb��.���Qp�-oA}�cXq-�������.x7�Q8N^����_���^��!�k,��#m(|{}e8'oЇ蓏s�#G�0R �_����C�6�¿�F}
��|�ͬ���k����c����S��_�������$�ɐ��ҿ����)���$�Ƀ�P(��a�<i,90,S�"l����4��Pf =���.�A:Ă��xS0�H�@����SF�eqE�,eI/���Ĥ�Oy����v�y�I�(�h�I���:�O�a�y�	Ry�1����4����Δ'?G���< ��������G>��ל����������������������%�9���2��?��6��YP �D <�A�]2�c�X��pF�(J)ϑt�,��F(u3��4x��PRW
�� y�[vW@Ck���~�jhX#�׌Ѯ���5�N:$�2:2�� �N�P>)�ҐխvP$�̗�C=�yrh��
 4��v�w)�����^��ޙ�n��g?��������s���~�����?���*A�!$����@����[��V�l!4�PQ0`�T:�F>���K���:�}��qQ�	�9�.� eWD�4m��ax$�~~ٽy����/�p�&vR>ʑ���d⧣��3�	�6D=x�0f�R�<a<@�Æ
���v���Eđ��'/�8�c�EJim�6�������������Z��9���7>�����/|�����Bq��#��u�o�fSf&doƒ	H'?��@ �Ȳ e��[����P?G�P��'˛��A~P�mu�+H'O�N��v��F��o:Qg�~��7@>���| o���øO��A�4�O���M�	H�,@~�D��Su�o��Nv>t���������6=���z��i^hh��εN������l�$k\�O�IǏ���fg^=�6֫����2[�X�"����w��TJ�M�m��PV ��aE@�:��t�
���r�(��mQ���]��3�ifr����@�:Q0h��@3�'�����`�,�1��C^�i�<o�h�j�Y:��Iu����>Ys^�;q�K+�ժ��xÍO��s�n#$A FA1�P �r���}y��P,�d�t�E;��tz^�#F��? H�����߼��a��#s /(�r��ߔ�6�`mSy�]�y����LN��w�C�q�8��;�emT��gk+2��`�t���N<�b�F���[��LxÍO�����HKkyOM�=�c0����CA~�z������7GҀA�q"x0 %(A���+7�����9y-� ����>|0�r�M�;�e�؉���X<��^-e1��/���J��G��L�_��@>I�-���>7 7N�����j=�����
�2Q O��;��3���L`�\So ��?�������۞{��ˠ�iP@�G㷃0�K�p2a�j�ŃnG�"�O�a��D��p�|�2�ax�%a!�Ep�a|��'&�i3��L����Y{���z���][;G�P�y�2��Z�����Mn�<>�a?�D�\�D#����S7�x�W?���;A^P�
���+�����킼�5?;�k=���	�y��g ��*K�yC@�d�C���=��cG����.��h�(��a�܉9t�H���u�Бk�}ilb��W �ʦ��P`�9��␧ފe#f�[��7���]�7��f��M���� }
����[<���n|�AڥR��׋pCȃ��	0�K��	��K�l�!�0���G��Mn�1�1gH���Ĉ��q���(�a��	���əi���^� yyD�A ���0�uo�СSpݍ#�14ʻA@��l�����O���Yȗ�7��>��w��J�X(�c�X�%�#��L\.�4ǀ��x|s�4<�
�-2���n���t��o��G�ڈ���L4x&cNe�k>[��o�*ɷ^դDm�8�@숾�λ�ayK3������ A��4f���l~�i�1�"��ȠCޠG�%�g�o��&yx��hה^*���rclLA��7������h����^��10���j��|�7�"/���n=���7�#���E®��8� G�OA^o[��(G;_{Mz���$&&������� //ʃ�Q/�-Ϲ��ق���`��V 
.{��|�τ�'����r�W,�)W�<&�*�2�7>@CBS�*N. `�0Lt~�-���:��x�A�na��@�Qax��(�� <�0��x>�/-��Q.��1R�(E��ȋgC��� 9���NG4�b��@��ʀ�=c1r�<�`�x;��y������; ��󾿙7�Ξ�� 7@H x$@��H�EJ�$Ǣ�*[v\��);�ĥ��T�$Rd�bI)KQ���-Y�e*&�� HP$� ����{�7����wg��r3Y|�ƛ�^�>���wt�����`GH�N������f� �稻�)<T�F�7���ٰ�|��S1��oM��Jf���i� 1��P�8������:E�2�칠��7��agNl��ɓ'S�f��ȇxHK~S�E��X�b�$?�#��)g�&�8�ƥ7��y:�����O.y��YzG�HԼ3|���A#m����d:���|��Ӡ_"RG-=��q����9�*'t
<�6�������L�ɳ���#�Z�R��z#�������z�V�4�c}+e�~ld���'.Y�f_���ɣǏ�t�{~�g��$e���������O�JD���'�۱m�7��� � (P���!gw������>9���'�$�u�8����.�XǄ�C<�Y��a?	�R�ӧw}��~��_س��T*��V]r@�ؓ�����e_�I�DrNE&m߃@�@H.�b>_Ȝ>s�d.�}����M7��ի�~�ҵ��x岇�[���%K[�h��s��~�NE"�Ql������\��l�;�өc�"҉�x�v�r?����M|����'����S�ţ�^{Gk�����˗<����w�ĝM,ݻD���7}�������*:Y�[FY]�ԃlo���l"KBR��4����������ct�B� �ʆ�u�.��%���U��-_��O`�0Ȫr�d��#��I���c==����u���^���ںz����ǚŨ�
���g8+��B�'�8�n�Oݹ��ܒ�|"}~W�؀�pKKH<���twy7�x�l�UC��w��-;���,X�OO�ުt���"�?Q彭Z49��S6v�HŹa��@D
�]��HAc������֬^s��v|��v<v�M�<�K���r$Noܸ���ۿ���[���yT��!I��x�H<7�1y0�tPy�*��9�8W~��K���c̌z�PP�t:SIf|~"QsM����L��D��=�O�zܲ`u��l~ċG6�t�B� �9���7��)���w����䦛��:��E+W��\�����y���._��x"�����T-/� �-�������h2 �K��6L����;'�x�c^�,��+���|v	�yh@�'�����;�6H�!iP�\c(�11T��Q��uT��ǫW�|�+�8f���7����k_Z�`�ߝ>��k��,�`�1l�UK9�& ]�!�ہ�@Y^��t,MT�n�����H>l?$_���^���U�f|*��r��A�Od�D��m<�M�i'7�����M���6�UnW����q�'O�a��rAW��֭[7m�9Z�jU����v'��	�}HXR�UӨa�H_T?��\B�N�.�8��"��a��qɇ�uD\���ʈ�7�҅ �Q�g{��ܩ"9F;r���F�9�mFš�P���84�������%�,9�➯W�mjoo<�z��ȹ9,���ӆH<�.N�w�>G�c���_΋�;�;��cI08��(��1��g|����g0@����l杋1���}�($�I��p;�k܋E�^}�Ψ\�#��|:�o,^��ŋ�1��@K�.M�_����K�ohH��2^�U�قo����E%��*K���A9�z�D-�F�H��|�r+��i�a�%rA(�NGjR��~��%�s1�lf]8��إ�9҄�x�~J ��  F?���#���w��N��s��̾E�����E�"��`>��a�5<T~L�ɝ�4_����Og&��|r8jR�ň��{�]�z)�*m�̿Nf��'ҷ���Gl;F���IF�$d����EY�:�_�t�ϻ���MbU�իWu�w�!�aSX\ ���y̼2� �t'��G��ؼ|���3˷2R��zN��!MR~f|�'ow����u���b��k4*;L��K>�7�y$��,��Y�����:.N{������uP���|�;�E���@9��Cuhb�6���-������F P�p�J�Hq�J�$T��{;�7@�\��9�'^7f?��f�4y��u���7$R*c�`
�����~�=[����o��H�w|���j����2�����~6��=�E">�F7�-��XM�װ���x=��d0��L�[r��:t(�O���dC�Ju�#�-�cs"��_N������y:<����#�&���%U@3>��p��v��0r�:?�ʁ��@�и���M��y���}�1�K��9s�����G�+�l�H_v_�ye^����WpB ey�]���Pӣ�%�y�l�cT�nQ�}��Bn��d����w��c�-m��Χ��W��K_ל��+����G k��ٌ?<8�g��W��E*ODR7�ƶ�,d@
2��}��ӡɝ�vd���4�.t\^��E�\((�y++Ԍ�O�G|e�#kĐ<��$���,�"�S�]�A�CH��!Ma�o��e�}�̆�����Hz�A��./�2Ij$�ޓR�a����,�|c��rH���:ruzkr��*L&�Kl=����._��7�2E"�P.d����֢�$��v�z��;1L|��l���PrirD�Df78b���4�ʞ���ά�z��U%�S��k���Z%�|��* d��7np2��7ӥ�AY�?9/]3 ��&�"��ӡj�U����Zڎ��A�oz��hH֏�g��0J�5=��U����U�����*{���@��!o�?���9������/�Kgwh��X����\�p�%�
x�P��=*��f|����K�t���Շ��ߴw�ުP�K�-:z��F�o�t8̰P���x�9^M���\�x��lޒ��*[V5#�S���1�3�<��MUķfT�,C�7�c'��3�F� :@x���;�wʨ:ō=vlы/�[*q�]�Ƨ�+ ��~�W�:_�L&͆�8N�>7��=G��xg����5)?�R3�Z.z~1S��K��in��h�Ө46�J0�V�	����$s��#G6<���?x��2ݯ�_>��^x�&I����:�͛�#u� �12�G�(�۲�rR.w|�����ɟ��-�P�T�!g|�1�h$"~�٥�\���V��L6�*KϥO���N�x�{�� g���'V�.[�]{�5���;����~��%znZv���?߱o߾�o���/_�fM�z|	�!O��, tj�ݥr ��
�4ƿ �g�9���4iF�'�����nT���ϫI�|� &���s���@8[�n5ߖݼys������{�_<���坾m��G��j��_nճ�#�{@dh�ϐ�^)�lH8�1�8׸�m��;g��������=���$�l� �d9r�	��+�z�re+-�&�*�:���Y'��!ɗ:�Gͧ�6�O$��{��{�ǣ-�/\u�䛿������s�������j�A�aI��]��W(�מ>ݻs��W���`�����6��n��7�~5��9w��p��ѹ�Q-r<���,���F��Lw᧍�w��$$�_���{��gnVeb�r�;)/
���*-28�a��)��w��=Sxo:s�y����fՋ$^~dd������ܹ�G����s��om�s4I�Å��N�I�k�T]�ɤ6���kv�޽@i�a&��Ӏ�"�P��)̘�侓v�;���Mđ?_�t�/����6G�w��K��=���?)޴샊���҇?���g����ǎ_��EP7b���z4������b��#�Ke3�۶lY'u�w�(������ Q`BR��Fݛ+�`�$��C�]944|�T�6u�mG�ݱw���ٳ罯�~p��t�ѣGH�&Odڌ#�E�lM�������mr�Y	7�&����Ym��9��O�(�j����ڵ�_�ԧ>5����R.�/��*5�ǀ���������U�p��h|$�� 8�z�Q �'�\�{����\��?�]�ݠ��FF��8p`��k�5��� %�+��ͬ
y>���Dޔ�w��j����b�,17�A3>5bQ�+��U�n���,�w|��Á�N�`�s���F� ױ{�^�]@IbE>Q�xwww���-L� ��w�y��v@� UI�\�rt]^�w���7&�>Cj0YL@��ԀE�ouur/�|�Ny�H ��X|�/�y^$j�88@G<�!%�X��
���I0v<pc��Y��N��X&O L|T��uG���
9^QN�"���oNC3>5D��U�6��J����.I�	��=r��#m����I$^__�w��!��"@X�n�y�b�ƍf?p248��9�hX�G�^}�Us���&D7�t�w�-��/�D@G Ӡ"��@�L�FG<��oډ�>��(�7���3>5R��ciI���>��Q�oC����I��֯���~�X���Ƥ�y��4�g�+��H�
9_�f>`D�j��e��k��v��iv;Eʱ9R��	�N�:�0Ӥ"��
S	��Wc�S�I�y��PG��7jx֏�֒�멗�k V;���7�]�L����<C<6*}BA8�����S�x_��W��~�oϞ��`K����6o���{K�,�k�����@�:H����k�뼛o�E�[%	8��>���}�{?`��N ؁̩4x�9eSse������Ͼ}⹳!0�C���k��:���(ͬ�"H�E���`�ۤi?X	=��Cm������������I�����@!��oH�[:���4�'�,�L&���A���xƑ{�5.G����j^mdgz$!�a�9��Eڌ�$�gP�8,H8�q{�1�l (�D�qyR� -Gܣ���L�T��&�������g_D
y+/Y��p�V��E}��[����W������g?�'����+1�1��aD���`�i�����0K �\ù��:&r$�k<�3�6&�}��.�r�#q(���8�d �8wyP��	�`x����Q����g��p�<��H�|�^��ȇ{�qyrteuq\���\�o<�8����}�ߖ-�K�/:��{ї�����֎.�w�Ĵ�ToJ�`p9&����'�@�h�q��9� �����>��|���V#]*��c�Kӕ��Hhw���b|��ǰ�|��#���)��[;H����@�`�\�ρ��x�q ��� 7xoM��p����������Vz����b�>��~}���D#Z����1\��FRH��T�(�?�aG��p��������mB�R��5�(ұp��s<��6o�|9+e�-��m���tAvݵ���[$ ��;w��]w���ޕWn��n���?����1W`l�7��<2 W�O����+�rq�^���]����)��q���Cv����U�b���y$Y߰w���?����o��HD3&�Ĩ��h*�ʅi��`�c,6�s�X�g��{��8:`r�3G������6��:K	���q��>yb��q����G��|�#��>�1��������߄����c&�J>��gL9Q�؍�I9]#S^ࢌ��)9�'�r�� A���4�x�M�o���P�/�+��aF$���G�~���^~y�V��Y���0�1�
�d��"y���eC��1�K�6t��M�������a�m����͝˦�I�A���v�hHRF+A  @E�&�x6@��r9��ĝSv6�;*s�8�?�����dlǳ�j;瀎�鯽�Z#��tk�n��Oh�Ȯ#��&gj�/���)j��Z%��,Y���I&�{V-Y���>����ҌH>5t �e����,�G�� 48L����@/���J�}�#�9G<�9�� 1�j۶m�V#m�u��wv���C�	���̌�1��|,��DA��?G�%"��8�sP�ݻw{�v�2y�,�.WWG��@�D�UK�I�)��3fȦB�͙��d�����8�#'�J�e���ӡ�$/���h�F3/"�zm,n�v��o0҅�ͽD<i�[[G�j��)���F�7sw!_��{�d��x�2�K6����������I`��`L��o���:/"p'%!G��0��'��T2���/��6�OI��bF�p�^F ����:(e��`�$n��2�T�2���l������/��{�q�~����=���?����/�����e�]������la4&�c ō���J��s� �ɼ�Q�) @��H($�N�+D3�v������?��^�M�����&1���i<#��o�2���Dr!�²����K����,h��� G� �P�LiI�K�=fV�p�3�0W�p_g���{]U�D����E�p/���4�|Q���>�@�|�rC��\^������0^|�E�p�u�o�*e޻w�w􍣦ϐ>�����H�����l�Yrx�RO���2�Ijw����:"���zժ�?��/֎�ݴi3)�)���k���j�s�\�������P��Ţ�O��Y�����E\�A>t�{��G���Gf|� Ml/fv�z^ ��3�O���h�A���f��j�T�%˽��I�a����/v�\��U���G�{;޳�[�r��]ʌK._�ԫo��^|�/���Řk֮2�H9`t4y��FN� �2��P���/��<�x /�fxS"�a�����%�s�O�	6��?z!�M���[F|?��4�^I]�x0f:)@���^M�8���_��Lz\G�������)��<HC?�9�,x饗��Cjj$.K�ٵ��$v&ia��&✵�n<��<0s�ԑ<݂V� �t��z�\\�D�x�9���#Rۥ� �S��аi�#�[i�"�t�hj������������7�q������Q?��#�K8L�wH����_��x�L�Ӏ�=�a.�w��9���4ŎT��=� x�ģ1 $�4�rp�������2d�3@�@�̼l�h̎'�)5�� �/���Vb^N �dp����q�N�3.P~����ϩ��1\w �|�@)�s�(�-��@�>>AN�P����BI������k�O~�=7���E�V��.�f|�g��k_��~1h�3p9��|N�Ø�(_�UH�$8�(�(4|Z��>g%&�b�Q�LZ��W�7	�HK�M�1�G#ɢF�!y���3X���/k��җg���q��uܕ����s�I`���L&g����$\'_��9���H\lL�uC>G�al?�K�:rN����L��pR��US��Z����[��ۻy�v	��NǢ�omݹ�3�N��$3�����������k��a�gz<�c1A4bߣD�Aa>�/����j�Tb���(G V��3��F�>`p h���i���aJ�5 �9d�x* A\��TP.�0��ە�P�Y1s�t�iऐ.����`ԓ#�9P!�LG
۵���Y)�s}���S�ԟ��>��sR�J=G�: �x�o�-7y6\~F���7��W����y�i����O~r��������� �0Ʃ]���8�nAh�j#��T�R�w�u�i<1�� �h��}<Ѱ6o�`���gL^���9��H�#�C"���� � }���cR ���x���VUy %�������Q&$`�v�&��>|ZiG����+W.7�S�|�;�3y3I�\��Lo�v}9y�G��$��%��6m���P����7}j������ߧ?��_��W�VRc^&�@�ƒ�s�*'�bh��y,�~����s�=:�L�a�
	FgRi#�h>����ۅ��ʃ9c�ej��N�X�dng��&��u���O�6��%M�fKc�$��<�h�x]B�R'P��c0@����"Y�<uu�o� (�N������:��:q8g��t٨ ~08�
F�S�o|��D�,A�:"Y�{)>ce҃o��*���c��������m��F��L�X����o��^z����0�}���ݻw�OL���9��Lo��H����x@�M���w�af>������w�kl!��QS�}�Hc J���O��h�@�QM��H�t�2��@@�ٳ�ip@u�̩��`g�k7l;��1� �g�5�8�l�;sz�1��$�RJ�:��S_R��	j�Ay>���&~.��o�$S�+�h��˽�a׮_�.���|��	+4��h�����ѳ������iSS���%����ȯ.^���/��i�糺eHLf� #ڨ��h&P�q�<�Q�	�C�nϋ{�W^�o�d@v��� N�QC4n)��(�3$u����@�.�nNq)+�?�/U: ;qhԄ��!5��*}T=�*�4��I����� Pc20|R���J
∐w������Q/-)�\l�{�P�u�z���S*�M�T.�� `�.�g\��8P���h�Ư��e��<�H$V��s3>G�qgeL3 �\���Ro�ˠ�M�a�����:�;#��/��dRc�H�Ӑ�����#��%i����琒 �����~�3�{Cz>�T�HI����݋���^B*�1=����!�8pG<G�N��)��R~:uÁ���3B�Q�Jl���%~:���Ư����⍬�����ͨ�#�� �	h*����6�SZ����xS��	�=�ޱ7O��ׇ���ߨ�@���`U;:*���%�hP@���"��d��*�$���%�L��>�������t <�z)Df.dJ����5lx� �lfl�c�/�EA�yhB��3I�Gd��������s��;y�W6�a��}�I�W5;��P>�M,w,���}_""�k�5(� ��B�z�_99Ra���O�v�����`<B�?�z��R����~��	d�f�9iC~�1~�&ĨT�<א�HI$,R�gS�� M����ᣦ<Hi�Əg 6�K��r�h�����~�<); �/8K�������6��}u���8���;]�fXu�=�1Ud��T� �ܹfT `3A�H�!p�M&�C4$�h���C���� 9�"�Ni�@F������5�7�G6��4��β�ä��� ء�w� (��.ã��9��Z$��Јʉ1��l�9��3�@����Tj�+o^�<��9ՇN������9���'��<O!�_�RU�"�WN���?u@qՠ�S���Y��) ��;�����k0 F*��J��?��X����ˣR��!J���q �q���G���H��wHزKbP'�	~s?�N�
���	)H>t���6vZ�H�4m��	��$M݈�}ҍJݓ׌箴��Ĥ�	ұGs0䮝�Jqt��'�f|b�Ķ��
�h��T�8�c4q $���~w��pL��1�&��^dՉCx���˦3����iD�9u�ţÒp1c��Q2�G�H��GBK��J/"�2f.�
�N��=���uI/��h���� jg:b���^2e5)l�Hz<��<���x�د�b���_T���^��6mG<�Ε_H�UH�v��1��9��T����E �|� *�I/BL`b��eO��Cz����4 �U�w�Α�ߦF�K^.p�ܨ�sf��6��%	iq�r8g�8�@BY �/6X:Ec��0��S}x� �K�Q?���/_�9�n�N�Ʒd܉gTm�Z�JB�3�S6.rDJs4�T�Ai;�v&]�ccD]M����@��r[ѵ��_�] !�0��*ȑs� 8w�9�w�c��%.y��6d�eb���(�` �a�Q�n�C6+ȃs��4��u�!Xu�����(}Җ5j�F�SePa vHR�t)�]Ulm1lM�	f\�l�z��ժ��Fz!��[|v�@١�_�Б�]C�\}X�C�&�u2�W�	�OӡEa������N��k3>1���b5_"��0��h,��5���8��#��1a<��\�����Xy�g̫����R/)�*O�I2CF�߇�|��S����s
�ϑ>�<�Z[����^w�<o^G�7n����c� �[X�b�#Rv�*σ�1�h���ލ[��n�z��庫����}�F���eRXv��y������Xl��"W���=3N\�h���#*�*�AE!��@Cܹ���d��xFsD�p��'J��b!�-_���r��j�����[�2}� ��4:�|D���d�!�vA��Xҥ�����+���~����[��w����9-�i�-5 cm!k'L'��G�ކ�H�(>�綷z�ٱ����1�w>~���Ȼ��[��4m���qN�)��Q�*)D�������%s�����u8�c�>�L�D\'0��ŧF�ۤ��
�8*M�H8'8�PyFr�"M��sNZ�a�o�2��X׭_����z��6���ۻ����Rw�
� ([�ĒG�e Y*i�<p\�sJ��uk����^������#޲�f�{�|����	��l	���X�+ݒ$FZ�c���՛7I�]�m����k��.Z`�&�0�=Oz�g��R���:8"�t���� ?9w��?C܋�c�X<�hK0�p�Qɧ�����x�w$� �]�i7��2&^�t˕r�N����6�-Z��m��ro��W�W�_��8"4j���9�g9�(�P�������-�VY�.�����yޜ�fy��n%�gȇNa�����O�+q���H]!�$���6�x��:��>�5�u�fkʪz�e5޷@X�Qn���0qʃ#W���n�d�F,���k|*56���B�`�pQq~�7�c�#���h�����$��A��~�J�Ʉ����%��jH�B�J~�]��*ϳ�,�͋AH������;=j'�l���Ƃ
ba*����"+O�ZP�����K�>�*/���Ǜ'�{o>�z��L�I�K�������(�y�c�H�o��2uE�s�����T6�6�)*���0*�L�P�X����i���2�0�
�f` �Ό��4���:$s�h%#�J&�^ϛǽ�o�F������q�Ō�7�<�y섗�X�S����I0p$_*Y|7���U���|V`R��L����;��=�:�ɇ4LGS��3�e}�eeP������{��� 8N <�nO�w��1����^��^/��zu<'�3$��&"�u-�N��$������p����1UUP}�c��\�OP�Km���Ţ�q6�K���L3>K�*�2ڪQkSX����ʥ����G빘l��� ��\�0��T���� �����>3�q��p*�:�C.SSvٮ�@C�v�L���-m���P9�3Fݹ�Z{��0L����P'��	�N�Ho:'�żt�sx�H��9��e�E8V���$	��Qc��u���	�*��_������s&����S�Y�Cc0u
�[�c���J���M�Q��)j�:Bg�E�q0�^��$�܅d]�̆���.3o�1�Ac�H�>�R���7Җt�v�=T�[.( j����Z@���8��ⱄ�
l�2s�Cހ~��%}�_�H{,=�� �=
��-yn�ǳ��PnV�p.��ۖ�@�)���P9$ʅ7�#t"��r�L��ۂ��Uy3�Ʊ�"�sۇ�XU�ÂX,�min9���t@Y|_��T"�2���(���v�I��0�߆��ƀ,-@`���`���0��}T�5�գ%��X ܈z��0�Xi2j�u��~*-t�$��,� ��=ǵ\I�y����\V��;&3�����bj���z�lu0I�(6�BL�0�N�^3��7��ܠ�1:V���t5ľ�ʯ�_����z���7׀!y�eu8�rD��x�K��(�,->�S�tF�$Wft4���A?���������4,>�$�#��������6��А8��R�\�niiy�����_/�olZvp�UY.� }�߼�_���8x��Uj|�0�Ӱ�����C��q������l�������$�Mި�&Lu!u�l��ݰu�idԖ��R}��{��}^J�ၺ�[��(�r��7�#�El�ʜ���^ /w�3�K��+�m�7O�x}����/P?�;�MhHr*gJN8�g���0~���
�!b����]ު���R�4���%���/������*�:Hj�ҥ=��������é�t 3����z4�GU�|*����;5W �m*�)�^�p�˗/y���+-��p!�΄�L���f���D���-��ߗ���U�7s� �Q�����4��:�㚓<�VǴRG��+7�~�?��n1���}�o�~�;�ެ^�%�f��<*lѢn��+7z�O�5�2u�#j�С#�(����L6xi�EY��kt�ҥovtt��3�t���k�?~`P��$��e�d����a̰! ��sRÃf]��D^?r�M-g���~}��������W^���G�r���M��u�/H[o��No��ETE�C�.�ۀ��=\.L��\  ��t�˷�r˷��ǲ��  4IDAT::Z���pNX+ȶ�%�1�������N��X�����MM�Yߟ��7oj�4� /�p��%p�v0&ӌ������+_��_��R��D%�!5(��h�Mh�y�OjBNSl�Ӛ�䒕����KW_}�+�h�����~�����;�T�CG�:�u��f� �S����V�CJ>�'�'	��ЪU��}������������g���?��'?j����mj0�;����ө�Ț5��Ɔd�i<�hԻ��2N���V.^����}���˗?��{���M7^��ҥ�v�>����~����?~������X</��/ė�X�_0oA� ?�o�H������~���A�،@�R]����7n���~�_n�z��*{�h�����|��駟�T�omkk+��m���6E� �IL�̞�ȗ�Xb_����{6o����_ޣ�?��3˾����|�?����n�̰�e~���UWmD�$� ^�Db)y�#INyg[Zچ�<��\������=߾��Y�vɛ���Z�СC�d2���ݻ�D����IU"~�U�s��@��-�����g������I�c�3s�d�ɫ7_�Ķ�m{�ŗ�m��ȮG�����{y��R�M1%#U���ȄXs�رUr:�dn��u��\w�Cr O$��B~h��>9:wN���u������i�Q�nҌ�z�Gd�F�?���s�?*:����$LQR�(��mۆ� ��ynz��'�?�Ѓ�O��
���2���A6�7ԝ�9~�����#����ڿd�ҧ�GF��������áP���ի�V�Xq��K/3�?��Ot�۷�-�)�7�4�3##�$���?sӳ�<��`./y��^w��ol�p�S͉���SZj=hi�O�_�e@���l���jo�����_�M>�̳�=�ē�F��J�S-���{>}��۟յ3���j�f|�4��D��ii��Mx�Tt(��:���z����Rkr�#�6o���;��Ayu��d����ʕ+/h������_���������̙�k�-2�����{��G?z���g�	�/���k��'?�l_o�FlaI����������ֽ������P�;M���������W�x�;v������tX�ď��h|�yN����GV���g���
<H�P<�e]a,���p($�+���P2�"�X,I$�~4���G���Gj����TI&�|.�
q5\4��d��s|��<s�Q�i�HT	g�����$�3����2��a��]��w"ǧej�f�򣣑\�OȖg�;,�@�$	�Ҏ<Ϗ�紴��~�mm��`�E݊)D9%��WD��X]���MeO�'�E�W+����'���=�[-�Q��ʥ�ҷ���
��*R�%ba��T\;�:�l�jcn3A�|�C�����p$�0�R��M��@��)�S_��I�%(!y�ъ�����
�S��<�<�z��3M�|~]]�H��L����
~��y�ڳ�=.�I��!�Ǵ�Q�n�(�NWeD�P3�x(i#�y�`�l�:����B>�c0�P$���[���F#�@bTG�N�C��?<<\�,��f���(��^1�My,i�]�}��
����f�z,ʃ,�yT[)ʴI�c5#k�$`��Q��F�i��	o��*.�LѬ_.�-�����	���E`��Y3+�*���=+%u���`KR�R�kxЬ��jN��5$� ���'` �0%�z�eXՙ�R9�,,�2�OeG���I�w�f�Fd����0�3xe��T܈����a.��҉��0X2��3��]zFm�Z�b��:-`�ӈ fDD�*� R�E��G�$3'U�ROi����Ǻ�i:�P�gGMV�J2�2�yǫJ�90���Պ	 �nm���M��Y>�����ʤ�x��P��+�w2�������`��MsD�Ir3�X�SkЬ_D�!_�V0a
�������*��))0�B,V��30���㬃(�kD
�(/�W�m8���E_�p�O�g����/902��o�a;���F�C8�x^��C�&��_T��D�Fͫ�%�ɗ����s�t��2�ER� �VE�a�I�R�����ڕ�6�:��D�`���|���%#ib�G�A��G��H>l=QN��M=J�j�f%��i����8gΜ�@8�bŊ�AD"Ey�|��|c�(�nWDr��!M�Q���n�Y�v�*�A�2g���UQ��p8�+��J7�P��G�$�T^^�6ӂ�}`ͮb�f�X�f�Xd��~
������p��+�v}y��x�Af3&p ��HJ9)͂�>����ە5�~g��c]/`)�y�zpp(�JשQ+nD��bT ����A�ޭ�tb����B�s��r|�DH>6�@�!=dě�jx� �mg�� �-(��tU�e��l��>�)��c5ۆ�P�Y�$�aW�l�o�(��6cx%�p ��lw����e_!�H�(��G�2���_ �
��f/�'��E�"�bvE�b��bQ�*f2�T:�p�U�
8X>%�gU��#�֨|.��Z!k#ü��p���Z���Bg�6��I�_��%�U!:M�'��[��E�WS
���D|�	�bq���X�y^��ds��*�v�kDcՙ�P�,����>��jzv�u�S�	x��NR��#��|��>��A�t
�peJq�����KI�wO���Z�]�4��W(,E2���b�6��`�-V }�e���l�*�#�t�K�B\"C��"�:��ZL�<�� �cg� v�p�Ng2�B!�f>U�@�N����0P^�]s4����Po��@��v���M;�hC��͢O�����l��|��g9H|V�� 6�k5;�6��'iQ��Ǭ��#���B(j�0�|�c�	͛��d]��P��b������}c�:��t��/z��Bj�b���S�k�{~�:+Ob�@�4ľ�|��3u��Ƙ>mڴ��݌�'���Sq�f�pց/����##���A�i�3��S`K���� ����I�V5�2$_N���0��:{�]�|�B|~6�Q0/��C^("�:�ܥ@��AN���g2	��|�D�FQ�|ؔ �1�R���Y>��H����2�V����iR8, ��/�o7_�9��U>+M�3�<������vk�b�|"e��&�x�B�W'U,A��p�ɵX�~��7��ď=Z>#�t�b�
tH?�����\�(%�lxp(4:<�g�qɕ���D�� �#�EVE5*pg����fqD�Ҭ_2\Whok���(�mo���)&�+����y��`��1Y��t��7-)��"���GbźX�J"f�f�F��b�A�|!T,� Wː�x'+_,��)5��[__�f��S�W'{5O�?���T&-�.�ݚ�|����K�1(�s̛��+&��E�~����P�j�)&�#&����dҩh&��8�RK�t`n����y��*�$�%��'ЙY� �Y)Be$�Ti�ޮl�T(��F2A��%�Oj�*���8�My^w�v�A<+�6[f?� �K�U�s�a9�)'kxC8d�I�&�:��0V�e�/�����6��)��s���9H�R�.VK�F0��a����H���oVJ>U�� ���1>Y^�L�il�E���}���)�D�J��c�^"��x�3A�|f�����oo�҈AP(�$�p:��H��3�W�]�- m$����y�m���ڣY���Ʉ�!u	��:���{���/��x�FKw+���h8W����!|o��Y>$�j-�1F�Ћ�HU�+�p��Q^i4+��ɤ���KQ*�8�O}�Y�tZ>���Eo�� &uv1i4ZZ�\�eO��3�#s��1ۯ���@IU�O���G�h�7؊�E�cs|�B�|>���� �UjLV�ŤK'�N�$M0����|���9�"�b{���X>����yE�� s��l2fFrx��P��k��(��L1�ͦ>���J�Ϋ�真��0���G�S�h<���n��:���X� �/��p�|�PV�z������R��H4*��� Te���)9:o^��u�ޠ�?#ۯjj�ݦY�px4KĎ455omm}����P,)ݮ�d�v/�����w-X����8)m^�����yj��m�z�οܱ�=_�|�U��>�L�v�Qͺ�ӥ]�vE_y��ա �*QW�(?w�^ٸe��R�����_�����{zN�:uꔌ����H�V�#l���}������ŭ[O��>d����:�A ����Q�̋��s�^:\�U�M�����E��esΌ�BWVx�"]�����/�Zձ����    IEND�B`�PK   J��XT��_�  K�  /   images/5be4124d-5fc7-4623-a6e3-e2055321e8cd.png 1@ο�PNG

   IHDR   �  �   �$   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx���%Yvv����ʴ�3=~v����X��p\��II�E(B�w�I���/P� 1DB4 `�Y`ͬ�===��?��^��1i^U�T�T�,�կ�|�7�=���9'w??~~|N�ω����v���~~|n�ω����v��_Ji����Q��O�������߳c�>��]}=����=��ۿ��5�1<�����˯��qЍ�����ko����#�A��?�~��-j����3I|�=�vnynoou�'�����+�^�2�m��cZ�<51O�eXS�Mz�-@��E��KM������S�������H���G)���ަ�$zu)�+���ӻ	w����E��ۙ�Wh�)�SN#
t
m�籅��-D�Ə1����c�2���ϣ@��(�)<�>���l2�*z�U]ǅk��~��;aT<������إy�����3E|��w.5��{o�M��T_�M�A�E�4n\S�i�����F�X6>�^��jʔ��t��[�|���kz�3�%&V���:�Z?�x�>-#��п��`.�kǝ��t�ϰYj"<�1�h�y��\�Y���lte�f��*���Ě�bI���*;Y�T�_,���>��G�޼��}�����?�G�6��w������Z��?$���6q;�M\��2&��,�9���_̃T�W�M���/��7�.D<�i_w)OR�7�>���}�`Jx��vJN�JM�� �~yT��o,���j�����������;w��:>w�#}n�o4��G��I�{���9|z�GN<��/f�.TX��R�_��Ny��v�$?$� ����'���wm��O�A�4$��;�
�	�4�Eu�XH�q��!��Ys���Z��zp��?�����������v�[nY�3�[�.���dޟ̫�9����8�OIu�x��1�x�ӌ+�.;v]����`N�v�`&��r�~~?6͹�X��߿��^�z�g� ?7�K�����՛eU�/uS�1)X7�3�&�&t��������o~�1�αM�r0�(�q~�:�~M&����k�a���_�;�7�~\���"��T�i���裏�Ս7����\��&������U��c�I�us�����ɯO�O�Γ�)����)��a�J~?~�>���)���K��h����Cmi����%�6��%�6�����+W�����\�oww��*�I��^ L0O2�0���~��lW'�p����X׉"��Z��^'d��}UW��ul�� ����J����)?�$�n�E���?/�k�h� ��p�Ţ����c��w>OW�gN|������_����Pxތ�b��q�pX��a�1�
�I��G1E����������'��g'�K�Tw��>kߋ��5:Vھ��Q�|��4�7��s������t|��q����W���	��[4-[�4'_{��[[���kD��3�_����&��ծ�穎ŋ�O�Pv�V�H�u����i���v��R�o�(���\B����e��S��Z��~�-�}��ݝ�7o���p|��G��ժZ�.M��h�΃�bM?�L�Yx�0�����$�dz��$K��^�k�}����j�;�i���}B��%�'������!�^��v���>�2"8?���i�S3�����r�ٹs?�S�>��3#>���Ç��HM�M��F"�kʒ'��@6�Qtaс�abNOWkR�hz��Ε�!�0$�l4r�X1�"�u��06_hjG� b4>�i���YyD1@x)�����U��T�~�1��‛�C���Q�sÍ)�ۼ���l�V� "�9J�Z�_o�e�cS��j����q���C������]�u��4�o�<5�-t�,�Kb�5���$��÷�q(��X�X���aDBj"ܺi�@0݃�MVMlvR�i<$Bۡ�&�I$>��_��y��u�޿H�msD�bN}�)	����m�'�lM��GtN��$�;�}���d���\���������g||&�����ǯU��eX`M]���x��ǝ��w�K^�#�3��2��])��)q�:��(')[���5�"���7��_���ɴ������q�j��݈��zcU5����u�|=6�/�}n�m�
��HֺpT!���4.�D`\��^|��fI�%(���r�t�^�~�p���H%�{�ҥ}��	����^MM�M��/��1��!�%���]��5�n+������Ȗ�v��R`���Q�3��sr��NU��!�~4�N�EV��t:-���=~���<���cz�.]������><�����𷖫���*}v���`l_���0b�Y�s�� ;��PW�_���MA�Z�W���lL��Co��E|dMW_�F���+��k�ԭlHhk.���_T7�u���k<8��+��Y�[t��HG�K��G"�~������w���A��Z������n�����b�G4"����u��Ms�:am�Q�����#�ч䘡џG#�nñ������� �>_�JL�����w�gt<w�Ͳ�H��%��1�+�J���N򇵿���� **��	��n�W����g�T�;�/�[�ۥK�������^����g���j���ߤg��l�wCW��w[����:�:n� ���zF�]M��rY��r��w���2������_'M���Gu=�x�|��k"�'u�i�NL���A���p�q]���4�p "�E��;綶�����ާ�}^����λ�}?��|qtx�6�o�!�Bul�v��k�*t�T��ڧW�b�A�����"��\�CnQ=�N3qn������vw������?|��Gj~�&�4�����灈t"F�G�k��~�\��OR��u��(8b�:�|����/���3
�_x���۷o�]���EY�7�6�0�kE+CϿn��}��^�l�y��ۿ�`3��&SLbSU���o��o�ψ�=7�{����|�+������RW��W%[r�Ím�1�G8�T�0���Ё0ݶ���+e]Y7�k�@�D���b�����]9�'�^|�㳜�_|�����	U��4�+d]o�,�����<�7����gO���_�����q�n4���r�F�)>�P��>_��$ݿ����~ϓ��"��H�~�t�l����v�P)>a{��]=|c�Y��O��gM���yoc���ln^xןq�w����X��-��8Ji���Ct\�q��sO$.{�'}.ĺf��{��֓��O�=��j��ͽ����I|;;;��z�Wǯ51�7�J�ԝ�֊Ǭ-����6���w�tAS�Y���Qm�]�/��8(����\>�gĥ��p��B�p5�5q��uQ�2�=W_�2�ț���a����������#�jN�#��U��-���m���?��Ӕ����W��9υ��"�Z.�7i�^6�cǩER7)8�j]���"�O����[�놜/A C�DᏳ��s1`�{���UUU��������q��{ظO�x'�uI ���ߘg�ԣ�_|w�{��m��3'>@����WSl~�&y{��8��l��@)��z@}��;Nlv��b6v�zT2�NiU䣇��t��NG�$�H�Ś���64"�zu�nH�����18�ܳ��oZ!Lq��kP����t���~�q���t�����9gJ|��a��keY�C�M/��>F|'�8�pP{�'�o0ɡ���c��Ō���m�<��%�=�c3�y�B&Z$�����#�!��}�c+��sN���Y��op�&�լ�_������7v�m��Nz�=��L�o>�_[������뺚Ş���Ҩ��F�,_׷fmg������c����M|\[�:O���˧��38���ʱ��¢���]��T�͎|M�6*p]T���3�7g�/Bܻ�D�U�ފ������%�~����wf�G4:8x�jS����v�UJxՇn#CL����V,�9Z��n�{�rݗ�;�_q_p�|T��'?�F,�=��#�A�N��sNyݴ:��O.������	�F��_k�}Rt��i^7�����z�x���{Ǚ���� E��~!s~� �E)�\B*L��J	%��ۋL�OR��;���YkɐĽ�HR.�;�?gr=пh�����Ń�j�㱿8�)�l�&����m����ΦFsy��!��[Pl#]�O0Hl�Z�j�镸�5E��<���_]6�7�Ų���ݣ�n�~�o���w&�G=��{��XD3��6��e��7��t+� � �����=M��E:dUo�}\���=�IF��9E/3��EH��Խ��3�๸Zp4��m�K$rs��VH:�p��t"g��}+���;w2GԳN�z�q���Ċ��*@���$؛����u���gB| �V��7SU15�HD^����]��2����"�ѷR��_�����+9
�{+�5��G��&'��2p�gU��[�|�>����^�O{�u��y��o�s�B��ʺ�Ta�!�����	�|&s��3)��K�hM6ZH�ꎩO�z̃�ۍ��!nT����Z,��`z�g�����s=>5���?~�Fݔ�G�y�����r��?<Lq���|憑@Zh�z�-�O|!r
���rAFu`�iLｶ��������=�z&�yu���̇�06��af��s�nB��?�����t�skܴ���t�����7�M717�3<>5���o���۴�_�q������z�I�+N����D��RN&��`P���oI�}-M	*�Y`B,������S[>��Ŭ�;Ғ���g�jXɾ�<Z����GI��=K�����~��j�w&��6�p4?�zV>�t�0�W����zM���ܙ~�ݻg����6�r��ֽ	���{��"�������O�߿��,s=>�ts��"��4�k��Ǝ㹞�C�1�����m���������z����8Y����\lL,��/�_�0~{:��g�Ν�����O��~kT@%�Ks�-�+wL�b~��6}�U�������L���͝`q�3�j��+�G�oL6&?�tFS���������oC1%]/7�O�՜�X���0A����g��$"���~f�D��b��3g����N����4�Sb��GS��i^j��>�>xtp�џlm}zX�����࣏��.˿�g�Ŧ*[�&se\nM-�1�w=u�k�ר����q���M�O����X� ��ܹi.��ߘo���X.^������������������x�od`2��Oq~b���$��,Pt'h�;?��qo"�w�����~&1�/��>�g�{�����_onn���۷o�����?<���t痳"��bj�d��Uu>i~���1��A�ωY�Z�B��.i��5�O�׍QT������w67���~��G�s�8�6U�f�\ϫe[id��J�>�۝r�7�u�Zw)tn��w�\-|=������5(��`�=+�-w5� +7"ݯQ4�(/h��ͺ�u���������}�gn�y���{:� �hs��{����yt��?����f�r�"1���<ط`Yp�>G;��#ٌ����"�=�kI�����Ȳ�'{�m����
����˲�����o�a�p{{�����OE|�L5��o7M���M�F���Фk~m��u�s��uC��`Gz1N2��:KS���ܡE�6cL-\��<ި	�&z���:��W��.ӳ|u2;�7�������77���S�y2v�����{����꣏�~����:88�ü/6)��"j�W]n��JG��s�>+�7��y�%���*]f@w���>��E�ln�����Wb"�0�[7�B]��\.�Ay��]�S�1~*�����|�(5�U,��k��8����\Ċ���j��v�5�'�&e�A#��`��w�TP_�luYh��פm�WG,����ܧ������b5�>O�q8���d<�����O����;��g1TU*��?�Q��W���ˇ��������~�6�E 4����\�H#7$�r�����I��D(B]�Pa�Z��g����C�7p�:7�s�#@;���dL���������>��?U��g&>�&q�W���2�y��~�����h�b7����Ƿ	n9�n^5�#�UK��[|!븪����"�s���\F艚�jua݅����w��ܽ�h����Q��$�����m5M:GD����(�<����)h@�L^P�\�&R�u�z�7*�����;���[�'�}�ap,v�{.��,�%(HQ���{}Y�~�h6{[��O�x~f�[����J���%ʛ:���c���k���])Jf�S]Ŋ�����A�œT�Ib,H!�,�b.�P�p?�"+L9!-~��{/�8��
G��fRmJ����Xp� \,H_�b�ج���${�&~�`��$�%�,<�4@�xթ��2��B�������T��2�6`�H[�(����ZK���Z��%�����I`��lD�yL[���kE^���x|���c�S�D|4�����[�	~qJ���ʜ	���3?����]���5(��5` �����r=��¢�Ɉ��rŁ�������颗Bĉ��2!j[Lm�����@�����l\~�&'���ҙU%1�0Vp؆�ԌH�4^��H�(W+7.rd�u����p5��.(��P��៰F'r§�iL�?��T����C0j��������������{d|���S�ğ�������k�د�`��(DFŏ:�Q�W��"��,YZ-4u�D'a��u��0��F|\j�,�y�"n�h�z&��a,�C��vqh��d6u�[�����eн�p���r�h9L��	���E)�"�Z��xc�mn�\1;��pfI��{U.���t�#�֘�o���r�k�_ǳtA�y2��s�d��ug���qf��7l��˚�q�#��7/�E]Uo,�����s���6��̑�g"��L�IO�5��K"2�5Y�yOl�[K�� �Uf $+���ߴg��P���j��N�GZĲ����b
��R��┓�[����S?s��ҥK|�&u�=��J�O[,�0�����u�0s�pT�9�Ͳ-����ϟc5�]N�l
l�|,��<փ�=��D���2ݐ9B"׍P4�t1���s�x�l�WU�)�9�U���v�36�Pߒgc�Q�B�e�v��/�����X.s�Z��6�]����<5�z����͘�WB�%|:�MB�&�D�+����&Ca��>��ҝ�oN������vP�®gJu`�X�пz����"n3q'����b	Ը�7n�)=�~/ž��%'��I!n��b����k7����,rKT��%?�s�:Ys��ٸp��{�75��`�k��C1�ʸ��D��dJD��.^t#�>bҐ=��̩�T�\dS;���5��|�� �H��1��w�D/|�n�գ��Ho}�ރ��L��S�����7{o�,��Z�i��`;�5��W�����+��S�eRj�FA��)&c&�բv��bI�Bu���>Y1b�l<%Sd,�X|y�%���(��d�,��MpWDV�X<[��c�O���	#"�UŁz��ZF���c�X�@��N�F����xg[�t�)[�rA�Sg�ۜ��6�Ѓ����L�/|n��U�J�k�띶��[UU�}��o��w�>�O:NM|$>f4/�M6�h�ٚam�6du�*�t����߆��l��Ik;���DHZ�E��>��| 8v�dāp���vy1�7�qx� "y1Hp�V��K��J�tj�Z��BD+��x2c�*UH3��A��J��ܰ8Ŧ'\-n~H:i�b�W��C����#�i��M�d3q��5ǥ���FθTj��K�p}�[1%��ahζ!��S�1���W�w#n�O�+����Ss�SM�F]��>�#c��}}��n��$}�����'�p-��)�W�B�����9�ʙg�$}(O5����� �E��h�=Lln��Y��rp�-�«ʕ:|��oEo��T�q8�Qe
T�t�u���Lgq ۗ�R��
��\O�q_�|�Ѧ��L,B'��ZnԉϞTY���I�هuf!�1 ��}�$�5Wi�~�t�����6yj���,�$=/��?�H!����<k�;���?L�d>(��O=C�3�DXDܣ�#�W�.hd7���	��?��#ΈP�g�Īk�)b�����e"��d�K�ש�:1��/��L� JT`h^-�7��p�<Q��g��suM�<��{�?�;G����l|27�U��4ĩ		9˹B���Hܢ?�up1��8����b��� ˫�֯/��v^pC�~��1Ϻ��@��Úu|M(�	��T��H�$�*�ml�`�-k��JO��FP����Q�o5j�;�/~��HW�QPƮ�)΍k�}�Z�Q��z���c��d�  ^\�8F2��mz�
v���uD���?�#(��O|����.����羭�B< �,ʋ-gG|8���	����
�OB^�@�RO`p)��@�Yf��D2'���'~��&pB��gE�G)C�D-��t��8 Bk�*)��C�ki���Y [�5��`l�"�Gy`}��\wF��*����L�(늸�����wըs�Ĥ�1r��5�d��������ݭ�����>������S���Mh,WIO�)��_�4e�D�J�X���g&����'�������I��'v�H���p�f�$�"YYt'IةS'v��n&Nh#x�	OꀉѢ%����ɸJ�`�UD�ә�#���M�muN�B@�x�pVKm��"��Y����S�vѴpY�������''��ԕ�~��uxbP���F�;NM|t�Q�%�W`�]�w�_�l�~�ayصl}������bp(p��I$cggǥ��m�Ƭ�-�K7��t+�tGs2DhC��F�0�Q��3�E�lwF+�j�G�n\d�K��AFH�V$zq.�=���L@`,Ʌ3���ə8�W�r�uv�9�?��W����X�Q1qK��IeX����[2�g^�U%h:D�Ɗeӻv]d��L���ܬ��$U}ݫQǁ��$c��j}�qZ�C��W�'Yz<mw����=aG�NT�o׷���*�V�_��{?fݼ�$�Q6��9��K��da̶y�8��G���i� =��N�����C���G�upbmR��*I4��p/)a�'W��͗w��m�?ě�	R�>~���>Be/�W}ú��Ɩ[���ZSw��7�O9�ZWW�	]�����P��s�u��i�k� �(�'�8��Y8�$a�=����N��Ϛ�w��<Ⱥ�6�֯�ǯ�3�N��t�1N|w�X��[��(cq��#W�+F.��Nc2�����p`�l\��n�pI��d�|�����y"-�4g��q�
�%��=�aG�sď�I�Ūd�e��J�/-���5r���9���a�F�'̻O4ޞt��	����u9�:�������%>O�,�cEO�'׺_�����$=��/|�;�a�(�Lfn:� �n#����ʜDnFę��\V/�b�r[�q#('2ߡ�d����!ȮzdUEW��$���p��zO�R��.�(~�Z�� �"�9��t�V�C��FN�]Țl�f�ՠ�qe����Q��Ӑ�|�dN���3�ށv#�9q>�A���֙���x<��$��~�!��w���u"�#�	*�ޒ8s&"��8�P~�s� I�,W��fL ⨎��käۿ��}Pk3r�mN׍9
by28A~���q�^ޏ=�R�|��\3d�.�+qf���3T�Ț��)iEWp	���Q�4q<�ad�#ڜ���y>#�!Ӱ����=��F:r�6�FJ��ppTJ�8ߺ���;�#���_��=��s\G�,����8�Ey�:Aw
��߽��=��wWo��-D�jY���%�F'�		�Q��xʮpP�,��@h�0LDs:q�2
�9*i{G��?������7_{ͽx�+H�c*�pH�'"���_��vǜ���I�U�?�>�ӏ��Ś�-H�9u��S=܈&�n��\9�ķ���q�x���#��k����'�8�d�A�A����X7"�ȅ�=�? ���{���MDw����ws�qiYt�$Q�I��u��}��b4f�	D(�C^¥��u.#x#'ә�?���~�T�w_��{���ŋ�cC=(��<a�.�V��0��m�5��D{��U��M�5�݈��B�1�E@�M�x�'>KW������?�-�L����a�+����j����.�şnm��|w�p��������݃���˯�B��rW��3����)
���T�He.$g�u���ge��z��c�L���Y�,�j⬤'^�r�M76�ݏ>f7\7_��?���ܶ ���9qM���Ij�gy�qX�4��Tǩ��s���Be��t77�A@������%��н��~���<��'A��h�7H!���+n1��3#��P�\������K����x�ݸ�����t�Z�e�>ы�r�U�D��M�/�WK��t���\�*����6YC�^�p��p��b�n.�F�ܹm���|���Cw�6IE��2=wΝ?��j�6�~nhAB�p�z�r:�y��B7�?���O<Z��e�}�މ��%>��P��|�����;�Y����o�G˦�\���Q����7���8�EO�-WG���ͷ~�-IB�}6�v׮�@:�����t�e���:�%#����W�W�_gN;*2�b	�=1�e��镫�YD2ƆE��\�K%�&�o����[o�%b���͈3_�{��A���Kƒı����)z[7�k���Y{w������N�j		�2u�=�ъi�i q}���Ϩiu�߭��H&dl QMQ-��/�a I6����EnX�P�9\%ζ6mPGh�b�9w�]{Sro�r��������)�R�c�qo_~A�t�J`΅��9�pקם{�u�6�k���e5�Z���n�ijA:�|u�OK}O>��ʧ">��j�"�9;{��^q^��7�{���0q�ˡ����z�[
ulD�*/<[�$W=~H��:��m�5g=�e,e�dqZ�J�]�i�.�qjeTw<Tbܾx���b7�HCo���p���:����SoN�)8��	ֲ�3w2s��7��/���O��Z��z�E�j���'�ly��N�P�e��軣��Z:,F!�$0�ឋɈ�_�a���f9��h�����8�/�mq��~���2���r��M1a"����o ��֜�i��9�*�T�ݦ���dt�'��3�*'�Wk.���|z]`�Z���yb��I�7_z�g�2З�L�]��A��Z���o1/�
A�I�_������qUV�ָ
p#�>_ci�b�c���nZ)�%q��-N�|�����s�d�����nqx�:+W͏�,n�K�A>d1�w��:��;��;󧱺�����pV��\?��?�Y��בk��쭾�1�b�s�#�e,TN�����&d"W\�����Վ?HQ�0-I:B���q���Z�҂��dޔ������4#N7��@xF�d�ǖ����ےNPجo�G7�:��Z�A���,h�O&�O)�}]zF
|�#+�eb/szƧ!_��U�a�����y���˒\���	C�qH,jiY|�5�n�Xuc[�_C�BȽ�]�W^"��>�^vB�6��6��� 	H@�1�y��t~Iτ'X�-P���u��N6�d6��3�N�_������\��j������!sќ���'��ǲ���7��ʻ
S��axN�<,OdpIs�gi$@��D�(����l��媃�J���^��ަ��������j7M�%�3gKA Y^<։�S(�<�g�I� �r	��YKC];�6��Xs��бx�e֟�~���I�Wib���E8���lVL���X�<�7F�㽟��R��zO;Wc�BUk�����L��愱�߅�뻊Y'�c� �)-��,�oVn��o�Ik���������O���<���1w����"��{�%���]���<C�Z���,B�Z�}b{����uԾK���3�_��!�������e>zs0Slu<�bm�\O�l��ec��+qx��b�2.%.�he�|�#�^9�޵S�s��d�G�{����\������զn�U�6������T�ϋ�;fI�u���a������c���%��?��#wb�,BY��$Cq�s���}�|��t�m�]���^�����0�K���]+�!��b��?�Ѫ!㺿�lq���G��χ1��~��~��������څ2����!t0���z�O�?	\6"����i���]%[��D��v fu�ƟHe+o��N��8�����t]�]�� b��s��U�T�(&I򉮫?s\�������7��̲h�d�U��s=�n8�v�dϩ筯�I�ѺN��]!!%b�He�9�qZ���*�'��������]#�7-��{�����N*D_�6��v���A�:��o�����?�u��#������s�{.����A�kH>)�i���97�]�%N6B�@�Gǻ��D0��띎N:֍���q'�����캨�w��Z@"b�yu/�0����D]�����z����9��/բ�gu��6H�F�l���-QdƊ����Uib��4dW綘�}���^��;��'��D1�z��d���>N{�I!M�J �sF�]W�[D對9&[6/��MU���*��؏]I����G]�c҃��q>�=�@��yp>0s�L��]\]��Џw�0P��7Qk�t!��k��$���{%��:XWڂ7W��S�H�kI=0�^Kx-GU����C�T��S׃~���'&��u�`��w�a�E�3�ZA�u��q;��{~�(D	�G�?���O�R���]��@%{^[�i�Z���r��\U(�>�9hk#�&�L}���X��A|4���w�o���C`��9�跶dQ:�߰�.W�QlK�umw����\�W�J:�\I&���_� �n6-�����œQ�"�wc�m@��J&�*�G;qժ&�+7Mm�G�\9�q�Is��< u�˥m[�`<�^���=���j�d�ǜǌӳ 5�~E�	��7��\�d[-�9b�O>�n�}!�̤眈����.�3�xh:�f�VҒn���}�zZ�bH�L�Cc��Qw��fB��%�o��\��lv�:��iR�L���׸U%�Ð1�<�w�?���8�� N�B�p�����������8�7�l�^�E�o�r�]�^����eH���>r���v�G���Ȼ�tɓE$��ecw��e�ҭ�hL#k� T�V%`q.	��(s�;���11�h!G�@�k&�B�#w��vW�]e4��"�fB���;Y�ކ�m����=~$��&�ߜ��^�bp��ȸ���9"��B�����N_���;::`�P�9q\K^
�G͑͜����«r��e��7b͈ A�O7h�N�Mz���kzFħ�}�4X/2_R �˅��jA������i��r���&�u`[�*�}�҂��FX(�<�^�I�<r/�z�%uj4S�t1�}aQ>�������Kw烟ЄG7ڤ{R�9� ���0Jxk�0�*F�Vc����ƽ��{�����u��cе�x�R ��I���t_�ů��_�Mg[46)�����#�}$..�7o۽������id"6���ڒu$b9�{��7ܵ�/r�S�Kz#x$������������4/)�{��6�TH�B�n�~nܸᶷ���ݻw�}�����`�ID�Be7ݘ�_|��p�m��q���d�+���0g$�Y���5�3�4�b�HaD<XUΉ�0X�(�����gx9v"���W�dv�rY�d�=j����J�	٨/��6�$�r��˸\`�у�ܝ��V�b=��T��&�{�/����଴�VKI���ݶ���&+x��so�}x�w���4��E\ �G�)�3�Q5a��"�)Z��zY�/Q�QER+���now��Ę����6HŅ(�H�v�&_#�B�k������	� ���G21�BG^��W_}�]�z�c����]&@c��D����̌)���,�K��b,���Dp��&�g!>	��A7���@j�a7����Ѿb\������6򌩣T��խbS3�R�	�?�����|A����g�Tߔ���61� ��������L8���k^�oNbv�<$}��M����N�Ѭ*%�A+h��S�L���3/�J��Y��ͣPd��D0PF�ʹ�Y��u������N��k)y $I��(]�F�,8&����w�� R"g��.Ȫ��<ƺ�9x�A�B��7��y�i��=b��G���O�4���!��>g�=�9�1�H]�1�P�q�F&�,��j�Kz��n��'�*Fe�b�a#�����������\��ۏ���N�p�����U*�:�B�}R�u���y�#kk�EȺ��[������'����Xe"�*�Q�-6����ߑ��UMbU��S��!�Fc�����L���X�s&z�QÃ�0�ge~�8b�̨������T��ZER#j�n�p��Q(X��|���l?� O�[���p�C��6�Ӧ���*��1���DY畬�r1��W@�H#7���3�k��ȳ!��h��R���;�;�~�F,U� b�/��u�ukqSx�a�ŀ�mJ���}U^�Ѱ���m��7c�4Hs+Y;����CzbC�^�ԩ�EyQF��nP�hb,����M/���F#��h�N��p�"�F.�L��ש�)�a%ϢD1,����������~|�~u�9��E)��l�]1��Δ��̼q`�0$!���4Ĩ����tax"�a�LWĚ�5�a�d(P��K�/��+��.~��FԢ��E�bW�9=���J�ўg]n(��>A�'�������B��Ud@.E$&�땤b��3��%ݐ��u�r|כ^E��%� ~�Ĭ��&u�Ri�8����DZfY�
��Յ��k��rZ�"jb��<N ��Y��I� jک���Z�7����P�bo�<N��9-3Z�*���6 >Y��W�I��Df�%qIwI�ϗ+)|�y�4��js���:�ωk���I���r��S	�n㞉 OC| �
�zhG����\�bƆ�yǛZ��M��P�3)����@���'�J�gҳ,�gܓ�i]kH������È'������1�T(WQj����ڂ�����"��(i� ��R�F�GB,pA��fX���9I���.q�&-�ǈ1&vC%�C1�Vl�ָ.s��v��Î����y(�=K��5RN��"�ȏA����j�g�9悢֍��_ 8'��ؙ���̦����wNfO��I�4��~I�F��|�߱��l[��U�z�(��5�{#j�(�qQ��>$�8j�5y�\"bb�&cU���f�4Ć#�c�C9\ �L���룶nJ׷1�gZW4���w� ��1�r#�}��IE�rS�c+R/F��Oo<�&0x?�(+R�H�����=��s��]N��c�v�8b]V3z��*�dځ��w8�&Mhf�R��?�a�޵ٔ�@����Þ@8.�K)��lbu��.���ͮ�\�)L�IX�ˉEM��{�݆��ıX���.X!G΁p���
9|Uܞ���V
1Y�G���_ �A�A|�Eɺ^5A҉�H�.�Bm(}e�^�\�:�Hb�X�r_iqQ�{A��u�M���t�-�P�ԕ��qm�'����Z0.<F��\>����Y��G�
H��Fb�^]I#�U��\	�o��E�e	�%�;l"��2���d���gU`������jD(6=�B^-k�$���L:��`����6fA���]\�ĵ1V@��տD�02qa�H:s�C�c�j��#����Z2��C�PѠi�Ub������H>+�1N\Qo��i	)E��9܎
p��U'�LaT�}& 
@���PZ�J����ڐ�G]�
���n��"��zNQ\�H��F�Y�%l_p=��Ok����Ym���(�]�pAt<p���y�.�"�%1���Tv�W ̅�D(�z�U#�@��ȹRO�d�f+�bkE%I�)���*6.�{����� ���H�f���!��X�N�q ��#>G��/�9�7�������GO�c��HD8��>m
w�֮A4�D"FmI2x�9k~튫�/�ĲU
��@�����?��Zq���ř�sL�&���5߶k̗?�m��y��_���o���P��.���b���(�r�W_�]�t�		�O�M�㦖����_�%w��Un�%~��������y2v��_cn��36�P���Z f��OZ����p�/_�5�nx~���q�nllʘirI�n���(U�0n��Kݗ������K������c�)~�J#A���Ġ�i�n�5W��j�䆮��������J��&>g�g�Y��J;j�Hל��]ߖ��e�>����}XQ0��xx�>p��l�	ӻ������{W�^uW�\��Y��0�e,�� �C��<H�����Z����%"<�`1T�㐾�A��J~�@�Y�eBl�r�`Oi�A���n��迶2,�%���!�q����1��&�3q�r+��x� �Ͷϝ�5�0cH],=�T�5Я�;wPC�z���o�
�h�0p&���g����q}��nJ�H��ZĚ)��z��'z�.�鄍Ɠ�|��V��A���Q ��E4�Hf/V�S�A��1��2����b���cU���韂$R7�<vX��:���d�|
]��(%�Z��7UhK�.9��~�tb\5�[6��[W�˒�?���`97�V�·.������p Z�IB�Y&;��
R*Dl3s�ĦK���ȁ  .,K ��"��b���sb�繩fgK|ta��C�G�B��7E��xH�'��DX�4�3#����B�[oز,��Q�!�n��|s� ��Yqlk�T��A��a	qI�ʠ�h+��' T�O����2�O�&s��>�&��鸶s��H8T��;��{C7\faF`��E\1��͌[<xu�H� �k��%�6a���'u���AeЏ@˒Q��y։1�c.�!�͉ � b}�v�]�W z��$�}�&K��Ԉ�����FV˘�5�kS�"|���Sα+9�Ƙ0	ⵓu#�<�,��Ȣ݋qo�+�Z���,4>��Zq��Hg�aQ�婚��[�����=t�̺�Hu(1:԰���H;
I���V�F� 9��2��W������J݃�Ym�G'"�l4�.�����w��++�X�Μ�-k3r�;6�!�x��U'�`L4�;�o�䳨]�mD��ֹ7�pWĝ�TV��A��gG|�5�l!E8� ����m'pu�6�|�>�Iu�%!�5�:��5wB�>ڄ9Z�UZ�9G�wi�X��δ�A�w�9w?WD�����|�	1�����o9�)�l��]�8k�\ �J� ��x�^pZj�C��C�q�E. Wݼ���U�V?1J�^��]��o��P��9�u�_l�	T
� 7V�\�ˠmݫ��v�6o�vJ�Q�NR��xAĲ��܈z���p����bft]����9�)��8�I���2�� �.�0�s-W%w:g�)�A���Gf D_+���n1�H�A��X}�e�E�J��lpF.�D���c.ͺ(��_Ծm�uq����Gc�9G�`n��.z��WsF��V��W5�Y1s�]{%L�(�v^̉쵬���dy��` �<��!ħ��p�����T^���;�o��9�p�>$�&��J��伂��i�Т5R018Ir��q�����F��i�{������'�&��TW�����|�r2\\��i��ba����e(�:%v��*�H-�8��,���6ٽ�Sv��MnK��ܖˑ4�02C9׫-/6J�����;��|�礛5���暺.a��>�]-@�|��YpwV�MPK��
�-�Э4y�����^rɠX�P�C�{�bB}WKr��za�XV��(9*�TM�Z����e�2#(�f�:�2+V�ui��5At@|�:��.��#���3MR�I[���t2�D�.(��R��;����R1�:��r�� t|�ԆУ#Y����D���NZ�q�~�Dx�1��`B��[c�Yw�=̐�۱ѣ�Kx���N�����S��	j�KdCEz�	���c�ܑyh@N�p$���0�^)�2ś����o�c��
�xwx�o��8���H&�-���h��:j��,�ei��U%TKϺV5$�]8�����"�qj7�t�Bβ�u�%xc�:*s�����e��v�$H#�rʆ��4=)�*��k#i��^O�I�x5Hp湓�BkT�F|�Se<���<�z�<S���k�]�����vx�y�jvO��%���C�!jY_�½�#t���#C3���=I�t�ʶc�lN�Kl�J�{<-+Vx4q���(��I-�,Krol�XW���i<IB��r�����xV�Ƀ&pIvg�9ͺ�I�%�%+�lK5��뭔U��\���$���S�v���fLi�Y��"�r(�����Vc،��֒��DF�\#�de�U}hR�c��![grdQ�π�M��X<�j��U�Q��,ė�����8G��%	�84�߉s"��9�^��</'��r�/l{��oP|���F'9!��o�j��X���s
R���1��։cH�ޑ�QsP�a�ԉn%Q_q���͉�r�}�B3�Z�ZT!�j���#>8�s���ԧ�v��#���t���c�чw��oLgn:�����PR3N����m����|�m�;�*�|݊fA��X��w�w�c��ooθW�(�w�'����������p9ݏF�F[������]�s��������$F)> ���h��8�l��^��{����d���U�EU���ƽ������?t��z �wH&*U�p�D>u/����t��]j�j-�`>H��h�v�{���6)oĎ'5��u�qpa�.�
��b��@�� ���"nUj8m�Ny~���'sfx:(�eU*Jz^<~��=x�1'��}N@λL5#՚ �i3=�����i|<f����o�/]8o�ֿԺr�"���K���w����sLo�X�zX�#Ttě�o��ɴ�	�Z���[�6�������/���B?b�]�������t��Mn��|�&/�3
a�-�[��Y�����������4g\k2waz�K�q���y��qY\��U%	�<��ގ���{��;ܠ�,���� ȼ�Xz�`�ELЗ�c�H�<�]�v�_�6ϵXN�)��U��WgM|���0��t�F&ĝ�t��;�9r7�%E��X_iX�b���Ieh�b�"�ȝ���$���?vSd��Eg֢󾍏�r�2Nt�]�\�{w?�����L�,W��r
�A+�\(������RO�x�!i�?qU�v�1�v����q�Wld,�����d���5���2Ă���X�M˜U*�{%����]2�8;��EB0�s��.��֔��u�	���"){;;n~��Ih�R�p ��I�dED��0�J�1��FO!�c��qJ�G�s�8�Ά��{��g�QN��l<i����ܗ�\�4잠D(0
�"#�w�̯����yQP�"j�������z�9�A4*�K4���ZX<^\ĜK����ſ,�Hvz��=�ySȿ�FE�2`a�:�Ug��[�%Q
�%�~�:�U�b���w��J�[n� �=`5��H2��g.�we�:�Ċ��
��p�>�aU�L�vj��^`	�TU�h+�Q���X ��|��.�r̜C}br���|N�/j�3��j!FN]\H�3p3.oR;u��P�]��J@X���!�Gsw4�g��r�$EjDY^+L�	1O
q3h��uԤh�؂4�@D����I!�FpI��ZQ=*f\M)���-Ѡo�6��p��b 'R ��:����驒�D���&����ld�
�0b� �1�;W���Gm!�L�� y暤e\�R���m/~�\7t�Z�zL*����`��@� w`]R@>y��3�|8�3�M7�L*�%��e���uI+8lА�w,v?��� }j1?t5�|x@ 2%�xQ�4JM�aUL���C_o����F'���#��tz�)n��Y��/$�?~���<z�R�D<tT����H���ر�bϗW��&'�!BɎ�q�j����$��Λ0d6�9�jbΑ�F��.�9�쵀��Zԭ�_��u�7�;��q,�
�qJu-�߀D�@�(��$�ٕ�yA��q���	rUA�΢�9!D_$�8`;�K�Q*V[��Zx<z�["c!�h$(&Eyi���J"!&ڰ#/UOMi�P\���/�$�Έ��{�iK�?�Zӓ�#}�Ƚ��w��G��A���t�.]��n�����*��͌�]H�	�O�8�D.�'��;��$_D66#2�4H�bK����_d!w������[�Cg���n�\��Z�W 	Q��J;D51�wU�y�N���T�wpp�sft���T�\Mu=dm@���;�*�K� �B'I'ס�Ȍ_��flmM�ܲV}2J��g��OPZ��$P!��w }��'9N���"�N߯�'ֲ8���Z���-P����4�����~�Y.�m�����~
�"�/R�}�GdIn��މ���Aۨ	��mNp�=mIrWR7K7-/4��=�pf�ݑƵ^�%D�uD1��Raٲ�BR�(i&�J��pl�I�83��:�^�9�81�@^��r>�H���&:�ظQ\Yj���tuT�DL�vWH�S�J=��R�a�ьw*��
�=Y�:uOY����9�q�B| �Z�W}Fzt�LCNHW<�#q�KK����t��Œ��o~q��h` Pâ�P�6/�!�b�VZ\_o���部�^�d��H�
y��<#)�S5+�c�IV8;'d��Я(�1Dz�y���y>��ܢ\0�ۜ�Y.�G �����xNA����L�� ���p�@6?�1��A��f��f.:!�߰/��B�Gm�P.�$N5$�.�,)�g��<z�r�g��j1��
�d�<�S%�$���D"A�'��e��.�8<���!�,4��RM��p3�hQyа��%+�X�?�;�w���j�.Nw����}!J��4�Őz���#Ql�"�Յ���꒳�h�D�0�(�i�;qt$��4��P�$
=x 48���b�cN:J\��ֲn#m�G	�d0���x�ሇ�ǆ�cX�m�[	��qG8�ߑ7��Ȓp].��>�}�ɳ��ܘN*��p]�ó">=���)� w�JA��jq��7cX=,:�doy׆������.�n�M�ݢ�fd
���3�,W���6
~)��%Mrqsڍ'x��3�@+����mďd6۔��	����p)9^`M©�K�t��y��җ�H�Jh-<���-w��5��}��E7����뺗�c�S���t�O����9
�-8�tŹ �q.��$���u�w஥tV
��3��h��9wp���L lk�s�Y�,:)a�����0kP���>uY�u\����sʄT�Cqȳ�LJ��[<�N$�|��[��|��A���N�z4�Blԋa�y���%�A�]$���ҭ�,j;QQ��
��z�os� ���Q0RI
�X�y^�\�\[��Y���P����ʃ��K��U��K/Jyu�J�>�U�޹Z� �+W���s�m�T^��j�i��q���kn�ſ��LK�5�q-!
�!�
������Q�z�9�ԯ���n����5%�Ə�Q̝a͓1�H�g��n���!�
gsDK���ԙc�P��]��"[�������R�	y�uw,�K+ ��V����SUĭ�� T\;q��i|y�P���ϳ>.��N?2�<�|��R0Ԓ]/���"�"��/�������������;��3I�V���/|g(q~����Eb5�/(��B���Xr�����R�T����͂�7C�ir6�������x��wk�j���;l�T�V����^גϏRB W�EG?�˜�%���<˓Cd2W�����ؕ\�_��n F��z��A������� �Ђ�����������`�\�)�����8���t������a��P�zX������-ū!�#ѐ��7���ε�2��p|��-,i���VL�L��}r���D`
T�6��k�*���D/��|"i�R��Ɣw�
{�-�9A��8�eDY�Ⲫ$[/�"�}�?X��F-����x�w͌P��P��y�d�s�1��q'��B��Ό7<\��n�9�$wd��⒕�e]MaH����]����кmFf5/��aNO�X�|w�Eږ����\h����(�MƆ���%�{����3�1�D��{���@���&W�ą��´_�{��^F%V���mi��F�JR�U��HN�1�g8N�E�gZ�x��f�&��	�:ײ�q���.�l2ϵL
V�{��(����g�`�ÎJ���E±x �*=��P�Lb�t�BZ�r�dpm{b�;��,��|�-�rf]'ڽ�{�JiM�"�%��C�0~��k�*x��<������`Tp�?��&1���a��,�����^���S�G�ϖ��8>8��dn����	�#jY��)�S�]^V)��[|CSta%�F�K-�о���\G��c�H9!�:I���졺h�M�2y. -(��k`���6��8�6�� ���W���cL�|U�Z�	.��`ɟ$
�kK,ĺ�� ��77t�%V}R�5���`C#���6'uA��eE��t��(5�(J`?��d� �[�Nu��·�(��4@�5���u��Z��D !�E��Z��#�MrjP�Sq>��Y�7�õ=C�k�!1R�
\ș��V\1i�;T�^6h��Z%x �%	y��P�FưxMRd�uJ/��~�?&p�ڤ�7�{u�Y���$�5��Q�ù���bw�&s&��sVܜ�-��K
��p��~�9�%�Yn���F��O�B��j��L3�d�F�W��(��i7?���ԝT�n�~~�w:�#�����[�������P1c��*Y"�SE�=�p#�[Vq ��]���poC��>���71	R@�f%�MxW.�G��ٽ�=C���7q�ͻ!����f:�~q����`/��L����#�p&�D���ja�n�$���mN����߀pf,��d�W,ciR�j�k��rN]\"ޙ��!��Bɒ��Z���I�Y[�=:BK^��u�|џ���Ɋ��Įo�>BM�{�LQV���ÕK��L6�����҉�Z�jՔl��9J�P5�Q�гI��0����V�i�����>d���{+���z�_N->N�IA����( i�g,�5��{�>�qOy-�;z暍rAAa睳�6|�tT��}���v�i7_���	e;:`�v�D�z��`���|�H��e��#\���6:[<_b8C�L���I�p�����T`cr�P��]�X"�X����1j ��3��<���qR�"f���&���p���g��@9�ح��?\=�,$��5#(!��O2��*��7j�����x�%�)�M�`����蠇"J��Z��ib%>����H�k�ьv�ç�P]�Z��`��Tn5���1�+f
g3X��xa�j�йøp�]K�|3�X�ln�"3��*w���$��!*�}yY2��e&9�qe�a�֢j��sc"0���n��,�dq�H�񌣫;b�6�E�nW�
��e�K���$�K*!�E|�$�B'%���	�!#�(� ��~Œ�%�e�5�A��=��9�2G�prb9:$MG�$��g��U[��3��p�Uj��ь���E�s�x\^$�,1�b��,�R�q�/Q���ʡo%����E��'c��)���u2��7]��nTK�BW�/�h�������ڽ���r�H���<"��gUA��gYJ�9,X�d
z0@��Q��\p*�@�*���Ð,��)^�h���z���ܾ��4z��O-�M���0?��p�ʩă9G���=D3�E@V0�`M#w�,Hdk9ȸE��Q���r��5��i��+�*�������
 Evx��M��p=���#rZ")P�ΒT�2.�y�ON�ܻ���|P�c��=���%�V)N&��hړ��Ͳҩ�d@���~\�uw��=n���x���hb�}9��G⍴@�� �����ZN&��_r���y�-�ӫ���K�w#���~��ݿq��yj�
��w��"5��P�����+�~����+\����"����� �����w�y��q�(�(�Z�D�{������N'�o��?vo}�+"v�S�bA�F|R�
�w��ΎCmjĜA�������l��0�nݺ��z�-������D���MR�|k�6����]��u�v��f��������k�$D?��&��@n�{s�`"��^W�3�o���p���j�	/ Fd^�h�i9w�������:�'�e�?�H���{�捗������~�~����w��(�[������:c�n^�ޖŰJ	@�p>?X���EiI���Dl;D�lƱ�N\hM�7���K�\�RY I١Ƃ�f�EqM ����>w�|���!r_aߨ͂6R|p�}x�cw�Ƌv����d��8��_fN�p{����6K��<�q���;K�#��>x�]�����y,BGc����ڥ��oI���\��5+I�B%�m����D��X�!E�Ro��r!9#���7�R��{4A�n�@Ƞ�p�$FAk����Y��]�*f�����I��d[��)�	%+֭�<��.�j����r����sn��o�5��O��;jc�[knmn�C�Mӕ$�ZP��D�Z�ل[�~���=�"\�{�%���c<"v��Iv�4/N�05Ё�NѲi���}x��������$�����{��u"ĥ��W~�]�~��;(!*J[s-�� [�*n�%�ݽ���Ã}"�'�c��Ľ>��G��8m�,jJ��`��	��%#퐸2�k�4a=x��,)�V/@W n�mħ92@�H#hI4��	��-rIʂ�;A\zj3$�{�S��S_J�t�QLS�[��8��N`RN���
Q�)Պ�rT��o�G����f���/^t��Dt'��(��"���΢R1"�+,����.q�w�����m��^�z�-h�٪���(��9E�����9oW�������Kߢ���7�n�����B���+׸+Q�F*�.��Ϫ���Eo�"�����I���}��I̾�"��A�`"Px矡����BQ�i�n9:gl	�e,�$��4m��r^4'�a�ꨒ<&�eQ@�!�,����b�UgJ|[[.�阮��=�tjÕ���wV���HQ/��{����}�[�r�G��n�kׯssggG0l��>����(E-~��kȊ�KYL�(����ͣEb��-�ė��U2N�0�b�����?�� ���Whg����5F�@����O��;����<_��ٹ�s�"�z�Z��Е��&q�k׮7�A��2�[F��W_��<��`��J�|h|�맺�2�&uk��J���9m�<h����DW���.����,h�;�����9S��i �೦q0X�.�+��b@����*�hE��������p��H���~��v���Hw���A�g�I�!��K~m������+r},�ڜ�*��C�3�G@J��@Vn�AL�����	aB���!�Ĺ����x<���H��v_��o����(�X�-�-�7���a�H�:ܹ��%��\��	�z����Rԏ�ƂT�B~G΁�vZ��I�T&Z׏u����S4�T�.G;2��+�:V���B��"ey��A��oE?�of�#<)pk�;N��ۙ�g0" &�������|��۷9֜5�i�<N��&ͽ��NϠ�EE���Y�\�u.�ϐC� 
3H A ��A�h��-�������GG�/��O?8:��}�pX��%�%YW%�gJ$H�$�PsU��߷��ggVPT�.�7"QU�y���^�֢g^r;�I^FK���R��*i���L/ �+�ɠի��T���n_s[ц�@��c)&�� �&��p~lD `I�D�F�(�����	M]�F����opCĔ׃!��C<��r�$�4X��5r�����n�[�Ꞁ�Uu��Q��P��;惭ӈN�`��,���7�DH|}�Q/N!9���*k��ܴ�xR�j���ò�/]Q�$�$���ׅ"�"t����N\,�3Ф(����,4�"�c��H�pŪ���5��T<ԅ�*���BAp��y	�Iī+=�D��/E�J���9�[2��I�v���Ggm�Ă*TxV��=��OV�� !�E� ����J�&�O������F-S'i0ڄ8EJ��Ԉq1�{�J�C|����?1	lDSJ���^!�Bl����v���_��$0����"�M��^�܆��
�	����+���cmZ�(�P 8��>�0CN�"ܠN$M87�������U�D�I�Cn��*S#� �F�7���ONK-@"������D���&V��_� h��,�;gC[1��ð���q.��!-pM\U��Ʊ��������)K�S��Ce�F�(�l ��.�@�7%	�k�g]�L:�eum����mj� �;�i*��p>(���%�+���k=>,u"φ���Rن�,���S��wg�<o(�ܝ�y���;����{���C��Io<����E�)'���=�2�V����~��o{"��2��B�G����l���EH�I��5����������oC���yt���Db�2�@<P&�Ɲ�6H�2,\�}��k����W)z�EoݾC�<�\#k^O�r�8���ӡQ%@]V���Vyް�H�rA>31�^EX�4��W�㍵VS�Eb�"OZj�XY�����zph�$I.mБ3�sͶ\ ZO�����T+�W�q%@�&�k��]�OW�U,
�`�s������?���x�[���Xk��Cp\K`8',]8bQ�bϞ=Bd���J���C��'N�o|����	�t�*	'���s��	�{�ؓ��*P!�T��.��>������ݹ=�+[�	���Β{���8y�bJ�e�M��g��qܩS�\��!�fx��UXT�M{��t�czޏ U}W7�+�P�^o��Y��d�%�4�Ԍ5�Vñ���]g!�[�K'7�9�3m40�U2)�ƚ=�^�iq�9_ξ�h�]5�S!2�!1;�
JC�q)�J�����������{��Y���	)��.�������)�N�+�=t���%.Q��9&9hO���9XZ6S�Οbn��C���Io6��[��FT0�_��ݙ3g��s�&���,u�{� b�!ϵQa�̸B"�a�ih�����{v�f�(!���p|"�S���.L�a�LoK�s^r`N�c��TڽREQ�6�YmP�j߭p�BuoE�4rE$)�0�Bc N����-�7�{���B*4x㛺cX���,�F'����Hu�=�w/=�"��b����db�Z*K�5B���8r�/���~7��+��/�dt����_�I�J=b�X@8�	Y\��2�{j��<[��?��Bط�@ �R/��cZɫvZܚH�������\M&�����$qV��60d�$��ɤ�'�q���ELP}���O���B�c���$ƞ�4MY
n1񴘧�V5 ��s5 y|	��>;H���d��SI5Z�]qi�Ub�P�B���j���"�d�dѼ�RClfp8�5���|�Bd��\�F�5Y����`e� ��\���DP���e04��ڏ��/��"�D`��sM<�����F >r�|J��-M<��R�.�Т�N�t��Q*��\��;�"���/[^[�6d��p�4R9D
�g���.4�7u�W��vI������*��R �^�����R�M�<�9�����9���"S�$e�r�8�JG <�&�ʭ�L�қ�<�}NT�4t�ma�P�G��}�.��M�q��X[w&��v�j]�A}�ö��A�JZ�6̗�+��6�R�Ы#F�GZKF�8�w>
��FǦ����iZw(�K�Y�
�/̾��qe
 y��S%Aobl��IKݼ�6L�Df���@����X�1�_�P��l��� @�R�M�o4���Ŏ	/vp�K�:A������� ��Zn�NU�uW�s��]��q٫�.8�B �A�)W�tIp~��`�َ�,��UP1b"�<k\O`J
�ן��R<��R[��n�u�8w���&���$�?�*7D�RI%�I�2No]�\h��MHH��bw�mal��.���ҬfϚ|m���R�;�i��e�H�a�Y<(��웑��VU��w�>��#*���D�?�f�Qw���J�^����X7H�Y��>�P
�m��{Yg��{҈H�zf��%eµ$v�4��e�ӱ�؋9rR�З5��ٸ�*�5�{��,�֊$�sc�5�S�S?׮���d�� @�8I{'�|��F�۷���+1P�#�P�-�'$Y�C�'SY���k��@�	(�� -ayZ�������� ��M���V�*X	5*%@A���N��;�3�I��2,HBa�xǉC)��i�JpN�LC�H�^V�+�:M$8��Қ:t�5�K�_n�Œh�����i
k�%&g͓�Y��MB�ăs���T�I
3FT�)ゟ�.�O����E�mw:���l���g�9q��!��%��
�:�� �P�J��.�Qf:Se�r5W3KϹ(�PVp�%R3J
��t�x��X>��i� S C��rR�D��DT*um,��ф�sj9�|W��Ҙ(�\I5�s[�";��&Ϯb��M��}2�'��6�!z_�' �o4&/�d��]�-f��:Ǽr����y��y�$Iv�YڥZ�|�t�^�n��礱Xe��<+�]Y,Q��>�� �ָ���A1U�w���;	ۉ�	tVC�L	�Z�l*1aӆ�m':[}�����D
��z|ZYȷO�.�jI�u?�抰��Uj��U��^�<��`��푔���4
�D�)7��Ia5 ~��*��W}"ڕ��`S���oT���vE	$�)���v�n�>@'=����Y�������p�,0H��|[���R�c!XxZ�L�3�(�o�x�
'-K%��^	-iU���Hˬ'�"�	��{���\]�fa�A������V�c*aX+ A�4n
���&�L����ĸm�TBzuA)ʘ�Q&�n�Ƙ����:��@B���f��j�%��l�Z��BO�Gw�hmb�5�V[b�˼  ���_����|��d�bJw�≶�D{h��D�k�f�Al��iXoڐ�p!�	��P��@�R���	���ګ�t ӻ߯��b�\�Y�n*�WL�l6Q)5s�Y�����I�@�r�է����t"'S�ED�Ot�F���;#��4�/��V[PN�j7���Rg��u�
%d^Z;�B+ T�d\�BE��Ck0Wڜ�1$���-�G����T�{F{�y�/�6P2YK�1`D_�ז�Ʀz����
�ū-�Wt��U��Obuy�-�͉�q��Z�ۈ���Kg#4��*�U�E"���w��$�Ύ5.&���
@��*w7�g�9�F2�|�J�j�+b�X�#�v���0ـc�qd�*��,/�����R���@J��= N�?���g�J]���e��>|��w��M.0 �7��ᾭ�����رc�!n̎HiM�eY[ˠ���Ub���f������"oka�羶t��͓��^��1���b�O�b�m!a|�ć�/MoY�v� 4�*(R'�:���nݺ�]�L(�T��婕?��녰{Eح��l��#�sV*����z����i�W�����?~��޾������\��tZ][#������oNTw��,d�5��ƻy��{�w܊�\N�Þfv���-O��nbr��Ɨ�"e��mFkr���M�����{��ܛo��|I�~Z�p�����~�p�;�~�7�A�z)��P�NHh7Ӎk7�N:�7?��HG���a���$�~�<���7��xf 0^ d^�������$���GL-���0]�������W��!�����
��D�iR�<qG�$�t�,��Ek��%�*Qenm�Պ9��8w�����5޶�<�e�5�I����g��{.�߭(�濢��� p�7�_s�?���Q��%W,��j���Eϝf��PrzS��&�H-% ���iqi�y��n��2O�g�"~7b�#Ԓ�z��(�(.5�$�0�=�zFp�o@��u�5O�b�f���A�nE]�,���o�ۙ ���kc���s�y�W6�-�u�@|���4�qaN]]-�HbPE(NC3����c����Չ(��t�$���~:qO���'$w*4��as�;�ҥK���u�qmĎ 8�:�AF� �KCwKs)H=YP�Swu������Uԃ�Db�n������S
z�`y��W��)�Ɛ۸�I�n
��sgVÎ	�aRš.�����f!�i����7@sJ*O�����	\��T�`�ᾄۊ>�6e}�n0~�����U���}�j�xP�Q2��o��Ћ��"k��;._ lGv�@����J/!ۡ�֠ǾL�Ӓ�P'��y�*��-����z���<!�&@�2�<��hCqmrj�0"l"o�C��js���L�St׬�P1/�Ҋ'��)nZ�삔D%k�}1Ŋ�,� �(IZ���\ <}�z,TX�I�âF���h�o�U>o�hH��I��'z�x�f�w��3�;�h�K� �p�AÝ�!m�qDh����I���ج�u�	p��� � {/��������a�D6��-���<P���T���Z���"~��I7�w�����c�O���2�~�����h�����@�N`�?�?�Q����Ϊ���	����L�n�ƥ�\��C�G��\�e�dáU���b	�0C�����k�����e�.g�Jf|��J�(n�Et|�k+qu�e��;�; �j�A�-�j�sR$a+��ei���	W�_��m'>N��/�k�1JH�K$s��	Z�[Jb�%]����괬$�Lb�֯�Zq�s2}f��V̪�5��Nv1��z',�Ȟn��"�V���{��1�L��s��$��3��"a��J�(�� M&�j=k`���u���r�-�/8��ƞ&ݞ�)�9�E"�e���M��>_i�7q'���+ij�3�a���Ăѥm$DWK��p 	4K�ɼ�����E�ܭ���-?�_��K���(�� ��j
�jh)1p
�����!^�6��Fx5��/���);�[ZXvs�g��{Cr�J�'C}�1�� � ���BU����P�d�տk�x�c�A�;mm7 �dy\M�D�q�Y��[,h��-�=���ޡK���["�g7�R�w$�r:.Ku���`�k�ڸ%�F]�:�Z�t�K�zͩ�'��b��\(���i.�;B|~�8Z*�ɪp���x�2]��RCQ���ؿTQW	��U�e��f>�g�H+����/P�Q�h|r�M����B�	vu��
eˊJ�I�'B�I;�ݵ��ʹ���HX�b���Ğv RX8�D_Y�@�v ��ǋ�<�1|����{k=��1�K�$D��S��J�4"B�>b,X�ӈ�V��\��+�C�PS���Q��`Ҏ���zl�1=A;ͣ�@UT;���'cB0�Z/�Z!đi��e!Lfj=k�U��a�O*��d�H�
�8,X;ƌW)j#����I~��6���i���C)�R�\�f@��k7�L���`MC�V�q�&���E.��a�2�w�Y�����:e�Vjh%F�O��"ӞU�CR{Z�Q�E���4�
ϠI��n�0 @�bG�ũ"H�n��.`���$����W10�PSԮ,��(�mw2WY�9_bQ�l_{�u��,�b��:D*ͧ��A��(��b;C��{�tc�~��z��X	�R����%��u��NW˻2ơ�u�:�����4������fI���ADؘ���D���~g/����B�LQ�'�VX�v�i��$�.9e!���PW V�:T��a��(��H��1�F sm�������8_G+Mu{�	�W֭I�}V�3c��0���������(3���\)ƙ���RUYzi�#�Gr����`�Q2�����g�+�G�����Z�&��z� :���K�˞�O�f��yΥ�Q��xSx�xS5Ӥ�|ȝ{���	�����a�m�tN�{��Q�qV�b�G%�u�ZYD�.�<r�4�MI��*�E�<�4���;��¶�}�eژmGp%�!O?�y79�j!�V0ବ΁�S8��8$O"	�E_)Z[���O��/�z���p�!�VC�قeы��y�*�� q9w����ԟ�!fd�lkR�Ӳ�%z���LqH�(ϝk��D�筽"*��Ô�7i�vQu ��T�D}4���1����IH���������:��~:p�U��M*�{��R���4#("��f��D��AˉG�2o�F/�-�!F�z���4yi)����敌�Ė��y���_���Y�� �C=9�D��"�8��I�}�X9#�A��Q\�%|��{���&uJn�,���..E"Y���qݞ�>`���`J��Ǧ��I�'�,��p%�!$��s�v�4��6	���?�T��%h�j�"�%�o���*�l�H8B��?��}Bl���f}�TEpi��ß.q�\�Ka#!���`e)t���$�����!�/9:���y��76����8�b�3�φ0�С�LUCם�S�ڕU���"���f^�^\e�o���^i>�z�A� �oH�Ɣ|E ������L
��-��F8���Z�m�mk��ܘ&�Y)�21?]�&r��LE�ğ�H$m���D,�N��w2qg���4ؕpTM�A�4�[5����r��î�$tY(�z�&҉"o�+l�MJ��	V�t<Cw�v���w��� ��Xmj�l���3�N �0l"E��j��\E.z^�]RjqM	���X7�K�{$�R{�����ڂ O5l���N x3U:I*b���$1[�D2�h|�Zѐ�Jtq@K|�\v��K��#F��%)FBH8\�����tKE�PAU����a�)�R5K�vU+2��p��i�^wj��مaQI�����Y5Uo��za���u}0�����F�D\��4J���i b	{��nt�A��s��"M��w����7C��� �Ep���bm�·��9KYm*=˞я䆜�΅�������8�պ3�
�MD�~(U8����t5,/VZ�F��e�ȷJ�Fȡ]���D]9$K�F��s�T��(<'$���8o�-V�fD�K�R�&(���3�?8\[:u������j��z� G��e�FbW�\����M�1��g%�>�,�*.�2	��)kh���C!�kJ�~?I�rg���e��
�-[�sRE�Ci�[�Ȇs*�팮?*J6.a9��BH�O��-�܆:yk��OU�Td�^'�833�V�*����^`UUP���ѻ/�̅B���	��(�1�J��a�kΪ��T�c԰zs��؏CcA'�����؇��K���V�Kr���v6˖�"=<���N�������cKu}��C{�,�Ǧ����#E ���&Š�u�n���:Z�����Fdi($	��I�̣���y�،�_�	"�ӯ�oR@Q��!Q��y��9�Ī�_c���ԔZts�S �ԓr���9��=I�A�O�&��3�t@�@�JWn1Z��\3��0u"�mQ������,TU�p�q1���:�"��-�a�[�n��Se(B_����ؒ�c�ė�Q��2�R��w�dl�t��n��6T�S�&r�=��AY s�J�>ٿ�#���R�#ʄ\K�Y���
;��%�+W`D��m��XL�/��J3�,�!��$y����M��8��j�l8E͸�(�a3IJ�j�e(Dɼ�OwS�+�P
u����B����u��r��P٪Rߠ9�i�:iȬeZڍ���l��G���,�aS��g��u��T�p�����Ȏ��DFr���n'b�����T�g3s�PlY���N��	W��~S�t8K8F�L��xɩHS�)k�L`�ε�T�& �����B����8�<C��hZ���&� #�"6��PIl�i�ZoY7c�d��W��?�i��ɞGb�ޏq;��,y��hZ�����6V���k]�̿j#߷<c)&N�C��N�M�e��N`l�.�yՁV���ًD8vXPj��)_�.`��}M*2�������d@*_�B��)*�-�,�.2�4T�K	�IߺBu��p�ܑ�J���~�J2�p,�>�*I��o��g�W��Uh��k�f�K�X��d��JY�$��Ad�2o�8`��j����2�Ӑ3��:(y��:�;MO3��HS٠��bE�۫"�J�� 1I�q8)��~�ؗ�G%��� ]�7�A�KL�]m�Y�Pz! �Dq�Q��ж4A��@xj�z�;+�U��{���V)aC�����~��>h*��e&-=�Q����_�O���\EQ��Q�,�$��W�j��>k�VW����ySN��}79��D.��zđ��IV&^�b�Zaz�FBrҁ�:O2.&�;�7�#6T��=�=�}�Ck%�,�AR������;2��ֺ�aN�Y��׉��,q�[�X���f��Ӳ�J���vV�B�pia���@��+ᵊ;�DE ���Z<�;D|inã~��C��Ƣ7��xӇ�u�o^��f*z�Re"����X)���9��I��g��j1�y3��l�O\�|�ݸv�E�)�S�5WJas�	ʊ=�Μ{��^�ܘ�[��v�!nɟ����p�ϟ��gǬ]��ΞuO?�4�-2]B���UQ..���f��r󳷙�C�'�����}�1���/*S��-\����R7��٧�Nڲ�A$��{U��L+�X��u������,���`׮]q�/}�^kPƑ�*���¬lDZ��H�w�>�*V���?xXbE:�z�M���c����+��_�[mq��5��,Q���	r�"GB\�Q�R:��=΅����7_c��L�%7�����^�;x��H��Z+kK�n�լ@��}��O^|���?����=zq8������K�@x�(��@�3�-Rd [d����k~S^'���UB���Q�X̵ʄ�T��K���-,���C�f�(��EM>��		��s�e�n;����uG �y��4��J�R���1rei����!�kIIVv��m�ҺՀ��/��n�Zt�%'���J��xu<��޺���v+�){!.	Hz�Nx���tKH(���\�R�
��f1#���ի������0��-��P�B��Ŵ�������<L1�M^nߺ���;�|,%�)
f�~�_-&�)�&G�����p+�K�ft��%�ih& ]DN�1�uʕ=� E�-.�����s^��5
�����f��.u}���P�C�E�hK����J}p�a��i�H*����Qt6��f�K��'%!���h�D'�O,�X�tZ�_}}���]������Иy̖+{�f�٥5��M\GE�X��D	�kv��nk(F��5e^�$��nu�	sJB����� vN,��80��A0��H�<���V���uIսy�,��L�ts��0�ؓV*���_�$_�Y=�R�<�1RC�}2y>���Bpsuႂ��(��Ui��6�)-�2A̩��P��`V@����e����F?Y����0M��GS�iS�C�J;9Ϛ����
��O'�$J�ۯ��,[��k}� (p�:���mD���C6A �~G+YɂV�]ZR����u�:2 *����Ї^�)׊T�.`�p$�b!�V@|�Q0h8����ie�ԍ��t��I�\o�}�cnii���B��Z�#��G����,��	��� �\],��YH�!�z���C*�JI��ķR;�鯆$,�0)�FHp����zx�D�	-�r�7\3kl��䦉ϫzy�ML����Qj�a��TFj0ȩ���>hְ =�VI"�ʾ�C'���(�� 3������pqsSKuNӇ�$��,e�2��I�h��'uWR�	�� X��{V]�A�����|���
[��D�?���e�t��d$��-�M��Ƽ~<����p{��\��fԚ�vpߴoJc?��c��.8����52Õ�L��\\F�,;	�YY6Q����kUx�.%@�K����j����A�.�A�~�s���(�`J���K��e�KӾ������J7��;+����7{}t���%��Ϩ[F�"}��e9�a:�KIu��Rs�RQ�R��&^%'X�]�c�3�!m�Kr4k^��e����?��T"��*zm���@�Й�>R4]+�`PY�	���� Ѫ��a:=Y%�ϴf�IK���%.�����i�HkX�͐�R�����Ma����$v�Z5�4X�Zaa�q�4�"�9���&ꇻ]�w��M4�� v�V��{�R��O�0��t�,����ĳ��]R,�"a*�������#��$�M��� ?]�TR?�G]��
@�=��
8S��ZrU�	�E�8*u"�� �Ŝb�����&yT&��
X��ʠ[��c�P�D*�b#�A�c�h��C'�'��P;��;��	뽎�kD�#oH�4�����##iڇqpJ�R���q���
���IH�>��9t{�[p�%� ᤢ��:��� ��dN��*%���X���B�-TܰN9(eȴ�O��9	NF�~b��|�Y+���@�V�o⧿���)��,}'�f�%� ��~��-�&Ao�z&kZ�DF�OdCkˈ��k���V�x��	a
.�a*���$��
?����־?5Jy ����ݓJ�@��� ����5e���E@��WO(Dz���
����3��#�����%�� Z����DY�!�N������
z�5�xcR�x�]e;�d.Xmܬ�RwWO�Lj���0��Sr)�D��3� ��BBO��
��N"ӂ{8�����!vP)j�,�ȯK�;��c{|J���7�]�-ѽF�Vx0'3���5��]�k�抺N�o��Qì/�S���b��F�lM�kF7R��,�fxB�k�b5W�j���9Ssa9��-#Y�e��*B��j���J�$*U��q��(5rk� �_��K�k�A�Uw[�g]Ʒ��*�FV2xL��o��_}(��Q�9���ysMb��7����VU��2��!|.8����V��g<QD�@R[l����lI
}V�����{AJ��M��9�C������v�K�$۫On6>���k��C��B�K	�5�ol���R\�I��Th�3,:rg��'幘����2P��Zf�6���5�+��Gˮ��;�cccfx�C�����,b��%��tMA����������6<��� h�k-�����%�x��6~�`ya4XZ���g�=1ɝ�������%:���.�W;]rP��yn�B���*�c���Um�b��?t�(��̄�Y�N8JƝ��������pc�>	�����	c�	w��SlV�&�K`]p�2nZJ��;#����C�K��T�Hi��kkB@�-������>��l�M���ּE{��9�����������r�4�~��jm�B�"r��ϱ�
w�|��i#�`���c�Wܣ��g��H�Hz��y��ט44�<����ˠM%d`��DP�%3�YJu�=3����C����H�<n���J��ꎇ�p�@ŷ�5B�\�f'O>�y,
A� k+4l�ԨI��_�U9��<V���&*������=��
�֎��v��}�Hd�9U�b�bٶ�I�U�T�$y�}��'7�O���10>
�/��`-G	���D�#G���`��Su�꾪��ih�*sZ?�y5���+kh�4ꈄǃ��g+�ˠ����T0�i�aUFsO�fx�8�ۈ�Ƃ����^ľS꾩��˖�Q�cu�%�G���R1 ��g�7W����Y�$�,�1b�B��cS��Ĕ­�t�\
d�����Y^Vzm�~�ߩ>5'����G�:�r����
�$fq��蝊l��Z$Ò0z>qVפ�����K��v������[[ʷ��R^�1��|�MI\��i[k���O��怆�T�wU�����vئ5�%5���A�~4P�Nm&~k>#wI�L$㭯����(9!Yf���n��f��V	�RDE֖$��i:5dKSm���`�ߚ�֥8/#N�����p�e�:��yN��«0l�b��ޜURtK�)�v�c3��FI�+�YU�;?v�>�*��t�;��J۬��9C����6o>@�$��v�?޽%Tb�n�~�{�rx���
�0�fzZ��Ke����ҹed &e$~m�$�)��=x'p��eVKy�LՎ^��>��A,&��2�g����y�iM�f{�LU���uN�f���IՄ�V�J3�j=X�,]�����qEMR��{���D�͟��H�s���"D��i������ȅ�@��!jX�[v]*��ª�SjcWDDg����kyUaI�u��<���AU�W����⁴{(��2�J��k$����I f��ؑ"��X�=xӋb�1���l7>���(R��٪��l�Z������:����D���1֬ѐ`q볫�-e��M������ݗ�n�'����*ݐ�ʨ���L�}�h� '�k�0���b�/�Q:F�����w)�I*F���S6���k��|�b��τ�mK��3X�sC�~� c)�w��5�IuLcđ�n�D�o-RxU�v�Y4�aM�\d�}�&�I��J��&�,�dz'S��F�]6�27���B��Z�@9\_ ��r��^��3A�>g��ITA�M��R����w�=�1�����A��$5(��CU�9�wD|c��v��r1��>���4�\B�õP�F�T�+#�@�:��s?��"�c�c��p�����ȑ8�]6�e�A���r<#�?�_"�٫*T��W=�z�u���T�T��	B{Ԡj�����bY
{v=�-�M��,�P�4�r����(�~=YI]�)�62�ߝ�.���-��Lf4�dZ��U�!g��K��]D�V���P8Xݕ>�z��:�}�1�;|�y����^g��h{3�i籹�i<Y��Gp֡�����VZF�έ?�&���3�ϹՑ��K��p�-����0�c�LFyԳ�߽��lf��!��<�-̬�M*���b�^UՖr7����Q�Z-�jX����E��v��E�`�0���v��n�7"���Q�5�HH2�a������<C�-�.���g�{ſ���FvO|��O��;A|ޒZa5���r�_��ET�?7�|UE���� GQ�Qܓ�&'�ry9]��2�.;;.3f?7
�ݍ��a-���q�9�r�S�M�|S~��a͔����7�k�܋�F�k��(�>s�����`jh����94щ��x7e��GY�w;�FL|�Dt?FU|q���m�sj���c�� �:��C� "y3ǎqw�϶r�Q��f�z�����Y06���K4`/Lq{_��;7�wk�u�&]���"������9q��TYܬ�1~��u�����5����s����6K<�bv����`�mb�����M���ǐ?l;w�f����Oӹ;|����׃n��"k��؆-�a:��6"���v��f�f��_�Q��Co��_�"k��r/u�5:�>��
|�Ǝ��M���bs+q��t#���k�ʰۮ��*ɿ���T���6G|�j�q����
'׊q�� J����fR[��������P�n�0���tȲ�l�u�3���<�k�Я�b��c3���bnh�꽖U��ʢm�r�c��emP�����z��|9:�'�f��F�Bp�h�i�F�E���ة�c��V7>DHT{�� �9���C���-W"��������\�����{�n�7��0�`�cs��\.��s)��jR�
w8�hC`����o�����Ԗ��ư7W���P�4�-�pV̩��m4j�1�u� ��N����zTQ����g���ؑ���ceY4�&.�w�ƨ���!C�=�ڻ��Y�Æ�g� ��a7A|�YUe�����u�����r�c>mBN��=�ݛ;��c�qO�[X��2�O���a:^�l#x�(bn�j���(�2|���Z������7��g#��	�'T���0��r�����JCZ_o3��s�X�k@'3z�mul�D*mO&i�%w��ͺL位|X�u�����e���ς:�	n��n�{j4m�1��d3���S����;�d�ٵ��&�����xr6v@���G��Q�O��ח5F-L��o�g�>>�n�ݽt�{�0�rp����yx�qwo?�[����d��,�����:v^m-�a����9����a�������UňՌQD����A��1��Qj�(�hԈ��\�8���m����
���Ɵ������D�o�ܣ����b|�Q�!�o7�K?d���or���6���[��RE����֭2�Mn8���!�G�����Ol����G-��u⅍w�FbsX���a�&��s�~F�w�{��m�I���|̨{_���݉*���z9lC�x���W&''���D��l�q�ɴ��~7��:�h��^��+���^�?��Ņ�s�ҧ6�%����7��0/����E}.ܨ1j#o���뽈�,e;���u_�������]'+4�u��:r�����������*k�jm�cE?��ws��wl�����7"�Q��6L����u��t4�����FcXǻ��h�K�FR��qӱ!���=����v���J�e��χ�M���a;N������3�<��t�=äI`6�PRv�R 1�����YO66M�>Æ��W�V d1Z%�����"۴Kw�<4HFs?� �6����������;�Fz��5�A�$t��kڮ4�O|��6X�4�a?ܪ��k�k���=�Kk*�o1�S�8�8�%M��Ȉ�mʊ��ψ�Z�#LS��u{��a�Faۓ�<���K�)�9/N�ح�^����b�ݸ�?��ރ��������Ū,�{�?��v���6�ݸF��5|c+�~�3۝� {G�b���th������ �b��1�V�Sn��155ſ�����v��}yy�Y��L[>�5�6�N�x6|��������"�>e :\�B#lKka����=�ms�6��s6�k��_u��XM���c��L:ȳ��y� �����޼iDh�k��F2�M�T6����]���ẻ��k����4����1?��;�c���7�&���o,&�_/b�H�tn���Z�l���l��ZFp�H#A�N��(�t[t�:��z��<�=���F�8g|��E�f|�n����)
ڵ�;]���}u�Y���6Zڠ�\8?"�����
KH����ǣ=9j���O����X���肰X�j��jb�n��agβ��hs*�����?���_<ןu�16e�z�q���W������5���	G=��_9�o�c2���/�l���IRwYg����x0v��wm�r�� �:p�@��f�K�.Y�N���R%E+��A�;�b�؄����O#.#,��������&>�i��=���te)-]'&�I��Ȳi�}�F�}��(�zE;�	a �'''�u�>���黶�k�z�/�u��5���"��&IЊ��wW����kmm�s
n�����%���ec������axx�?Ȝ�-���V�=������Ӵ�(�Ƅ�}~&���I/J����Y�����N��A��hPe���h���y�ꫯ�_|� �����;đ���ݼy�nbBy��7�믿�	�җ��;���쬻z�*ϳwό;{��{�7���B˃�_�[�o]ciqE��~��izz���W��=�V;h���=�Æ�|���3=�{�9���<�������~�~�_����̹�����$�k׮�wϿ�>����x=��#$Z,<�:��?�y��/<���F/^���9PW !��y뭷<wwG�QQ[E�T6xm�%N���&�t�{饟���{�:|�?~�}g�����9��˭��mw�cK~�Dz?-��n:���w��i��I6VU���@N��8�?{���~^����:czȿ�*�q�q�zL�&b2�H�=�������Rt*�p��@l�^�\w�̺7�x�=���Ȇ�0��+%��3����GN<L"直�y�&�o��x��o�k^��anX6 b��������/=�M�����*�;��7��w�n�p~���%��g��z�a^��?�w����GQ��}����_z�.'AB��<LMMs���\��N�:Ź�u�;x� �su�{�ݸq�_�!ε R/��6�E�5���я~����q>|�=���_x�K����@�e�U�&PX����6����Wl�|�'�M/.����ys��m��׿��w�q�����az
�_�*'����>���ԯڢ0/,̻��׿��qv��|��c�K<�x�	� m6F�����������]��3��5�Ϗ{ !�(��X8K�l(�Ť��b0�\n~q�MML�۷os��,�<�~���ک�����N�8N�ѥ����t�z�/�������Ƚ�^���{�x��Ӝ�"�.���v;�f)�@����}J�=���7��>>{��7��]��*ظ�h�Sq�W�^vo����ȯ�Ν;�����tٿ����
��x`��� �����Fu�׫�ꬭ���.���[�ka!���5�|aa�����~�����u ������ q��L+�]Y^�Baa1�gΜ��%��a�Ο?OB�y�5 r��������������݁C�9��#���?rO>�$u�K�0'�^x��C4 �����!*q��k>Ä'^�J�����kw�pB��[�����@_Z	������{��������w��F������ַ��^��k�H�H<'�Otф�����=���r�0�-7w;J|���ʥ�_~��/�'�Wd��]������7~�7��ӧ9�?��O8A��=É�v�*'���AGD7�eOhh�����Z��I~�{~�/yqw��-���������~��5�8�"�| �`\Dx��aqn�M���̦��o�"aaQ�끋���?u�7�4�.igc�&��$�w�y�^D�����pU��O�޺��a��[~M��=�>p^�8<gO8c�����������ʹ�94�����h4����83���Pgo����	U����8!����+γ�\q�.��߯2���%>?����zz���<�a��s��N�8������[��[��炓��Ʌ~����V�/^&Q������9��4+�3�J��<У�>�� ��	p.s��ĺo�\ &h����w��@�{=qcAh 8p�cG���8���y����q���t <Z����{��?�)��ujraXҏ?�x�l x���G�`H@�y��<!���'����ȏ�Z\\v��u�,oǺ�N���i�'>?�����~��_�H���LxpX�{ 4p$,&�� r᜝����CĂX>���Å�s\a}o��g���"@�7��^{�5�a��a��(�w�
@��hC��=��(�8E�Z��:����+��B�����O]��_��zҋ�cn�n	q/NvG����	��Y!UE���7��R\rzj�{��繁
uЃ�aca~���\���µA�����5���ԌWc���Ȟ�=r��} ��ް�C��{Bj���'�Nr!,>�������׿�E�C$�T,�?��B�H <�|�p(��j�6�ׂ�FX�%��<�_�b�+I�m��s��Inp-�����.	 ����J�����7>�q3���^x��������'��Ïxb~˽���\xl0p�\}�x����A� p�D+�&��~�=���<��������7���� ��h�p�X��\�>� ��\8�z����:<:�8�y�A3��/jj~9L��U�`ך�'=,X���qhJ�7=g��ߛ�����|p&�#�;�&[$��*9�c�=���'N�t]O`�x��Ƣ⾾����zkt�sͩ�3na���ځ,�j%�`,��ظ{��w��>�u����A ��� Fp�;�`�>�=� +�; �Vk�:�D�����]�|�=������ܻ�'ב�ܭ��|}��Eu�g�x�~%��\ԴY������˹�����=����/��H�L��XS��e,��ϰ 𛁻cQ�x�P��ۀ���	g-\��<�м���9�I����Q4v�u07Qn�����=n��� ��j��T�brl�E�_ZX��O?�$���E\zff?}�����<�'r8�9��C!����B�ȝ�7Gn�k�������b�%10�f�'�	pB��f�5�U�	�<o��l| :p�����O�%�(��3+��`aaX�ىI:q�_�}�q
knϞ�\DL�/~�����>	V��1��~�B��Nǵ���u����2<�	�D�a >Z� 6��+<�2�����e����2����c��A����3���y���=O��Ǘ�찰1�;�{��W� gZ]�;�t���nR�߾}�	�C�}��.P=���2+��:$�<�9�1b���:>o��#��?��{�r��
��]�W	��E���{�K��z�}a����z���w�>/�$,�c����H7�$	�D��`�a0h�p�~�?!.�\�D.��.	��s�D(;uM���|uK����qյ��F$Ĵ�$��` ;~�A�{�oem�`�8m�ɩqw��6��k�ۇ����p�x��O~��;;;�g������U�/�̸6�qX�àњ�\ �L����t�����;�Rb�L��h��80�I��������$�[�s#`ῃ?�&ـX@�_b�O��hOtND9`͚�����|�;:��Ϟy\ľ�����Н,�l��={�H�Pp,˂��a,���>�>�ē�~���ݜ݈ʈa�F"�Q���SO(�=1Cl㙠��{ �����-��������y��� ;Ǯ��2��7�f��L�������4\-x�5��Y\�v;8��'��1��k�I�~�������n���k_��NL��pn�ۂ�ׂ��5Y�yN���s�=����>�>3����0ݏ���qb����lWǦ��n�*�g XC���� ��}1\�ī��s�P#�l�9�߁���O_�~�́o~Ӓ�#���ź���w�����2?q���:+�t7�W^�u9O��k_���������WVū��	�k��81� �q��ښ���2��By��=�2,�m�c�a"�D:�o��Pp��]�qo��N����S4c ���Z&��g0b7�"�cn&�FXD�4�w�Ǿ������y�������:t=��f��?(-|�����`�z��o�(���؎��a�"C��0k�Fg�jgz��6>�a�	��A̾�v��s7X4�J��7^���w�x�����h6P)6]�k���z't4<ϳ�69�����c�ⵕPť3>p�a��Z$%Fw�C�Ҍ3���[tH�b|������^�h4`c�;�^x�E���*l��l6i��3��\ 6S�Al!����㻶x��W�U?�qUµ�	M �*�8ވ��~{n>"����lC�ˤ���C�&s��؈saE�l�l�Pذ�I�*ǰ�\�~R�����:e蝧��"��柙����g|���juK?1+�[DC���_����7�I�9��\�V��Fq��-"�Õ�08ɮ
���D�02�l�m�#�r�bUu:#�@<U�P�^����U�����ńi	JvO�c�	ۤ�����8��5�
�����S*�r qq6����&�����ϋ6�|��*􊵪z�2��p4��O,F����J�r�_�����ZI8~�z��
|b(�P�u�qS���p[�hX�FXX�X�4����8�����3�l��t#�8S/F�v>���t0d E1��p��sFb��4O钵V�$)/q�;��WWw����@$�#� ��u�f��ϓJr20%y&�g"7�n\Ot8�)@��4�5c*F�>0+���e��OO�yf�}���)�p,&jb�r90�ݓ$U/��A��9�ݣ=ð�Þ��m絍a�/x�g�d��:��%)F��9,�kV������v���W��;�ؾ���PKw<6R�~D.�>�cg�ʘ�`�3����̹a"�A��I VR�fM'6�ŢMN6֐���̠!1���kz��D@+t�Kw�pB�j@�˞�dt�9�ca���b}�Dn�[��#Z޴�p���:emX�9 سg�;>�ˈ�+�^���4�=i�W�����=��6���$A��r��I���\�g� �7��8�5'7 Vc抁�
aA8�a���.т�Qd�����m��Rl��E�9-b���՛[*�>j��pSۈ�=�k܏�t�qg��Į�`���ʄ_��%v��xq�^Cp:��oi�WT�9|/"�{����A�<>�΁�d� hȴ���� �?8��3�Neć�-5�h;�(����<	�Wo��T�X���Ng��g!>���=��{�f0�e%Ǘ��s8p�>���^uO%k+kM�[��O���RdY�ʧ���������D%~k� �6���D�����65F�3!�fE� J��5>F���beqi@d�:��<l��Xg�fg6P�����b��nP�AD���O�������jlw�ݯ}�k����A�I)�aDW
lG���J� a%��xl �����
F�f��� R�|��1�o���E��  �3"�/�g�d|%m��y���f�G^4����M䎪�0<��Ϭ]�E	t�7�	���kk�0�r�4��L�i5[��S�Q_�p>�A��U�̻�v���� �ٟ�E?M�n����njT2�A��B�8@t���	�c���(��� T�'0�D	"�[[^[.��x������m�j滼W�~��� f	����T�?S��v��"U�R��;���ܲj��<�w���"����=�6�n������>U����h��P�j4	����!�onp������A�[��&-��]S� b34�LN�q�Yzq a �oa4�A�?��Ȉ�k/q���11��-��>-���o�����"���|�k�Do 'U���.T���n��#�/�z�'�r[�h�;+�>Uxy�4��Z�&E-�X�yR�j7E��~���>��7o����)<6=������L��@8!������S��(gQ� G�#�HF����6��V,�aUE��8~�����9�06�y B�հֺ��]��h�cbV�oN�}:���6����k�2|a��ٔ�*a?.�XK�� 5�
�����;{�1�O�M@ o���5�O�:��o��zэKW.߹}g��}�������<�n�sv�96���I��/9Լ���s�0�mA�q'�f,���B�����4��ㆵh)�gז��"�.�)�*͒<]]Mw�����jY?�i>4J7|�`�xQR��Pq��P2��x <
t4p�n�ߙ���Ut{LMO������䅃-f�y�rg�5;{{���3�ss'._�詥�3�/_>���rȋ�	,"��<��C�@ 
ax�Z�I)(�;����6"�������r8$��&�b���<M;��χ�u��/x���_��0�c��$*߄������Ð1�J�"l��]{ff�O=y��Ν{��ӧ��*����Zy~i܋�����_����ݻ���녏��: B��:�B�|����e�w̵6�p^?�6��i����3�!3ڤziUzyR�|W�݆�E颱s/Z�K���^Ԛ��2�`8�ګ��5�`nz��ˏ�oO�x��O>y��0�E����5{���k3SS�O�|�g�����	�w<Ab]�V��)�����#������2dx�T�B�|eUfkk��G|Y�]y�'�^2ʚ��mv+ͩ�%����]2�U��Y���rx��ز'�7>��9s�����/|��V���0;?:����O�Ͽ�n:?��{���������Q�{���Y��mڔ��\G-d��|��|h���j�` s��w��vp��h�>�-7��-8�����_��N��DPy�t�ĩS�y��3/<��S["�x�9z��;���������?~䣏?~���l�0{�7��w����A������N2�~\u>�<�u���'Uη���S!�"wH|��vGq��ߣ{k��u�b}��so}�߻��n@���2���~Q�>{���:��?>���Mx6Ν;w륗^��^��7j�y{��k���K�_헓� qlR��	V�2�H��]sX	��0̢,w)��Ȏ�/6R��m�n߁�q�7l�ˆI�.>z�Ξ=���J�q��ԕǟ|�[W�^~viqq��cVm\���x,�#���a��L�w����~C����u$���*O|�	�`|jbWFzLH�;%9M;��5R14b�d~.��lQ�f�p�`X�9f�8��_ċ'}��'N�ٮg?u���O��>���_|��{��3�����w��(9)׵!����u��bo�2�܃���2h�Zf�� ��W�D�cE�^��y�w��-�,ɢ���ۡd��|P\1��jeb�/�n��H<G���减?��[n��'�[��x�_/}���<�;���H6��R�0]c�=�8���A��G�,��|��ؕ��Oj�Km�u�x L`��>�&�4�l��4�g�̪�e��ϋ��ӧN��ȑ#sn���?���o���r������Y���J�Y�n\�b{� �ü�4ߐB�N�@���>'3j�e�j����@��0pR��岦�hLGV/����bnn~���#W�N8ҟ��cfff��ѣ��sv��;�����Ct�\0;3��v�n���fi�#�%%CȻ����(�&:)k��C}��^�J	u�
����z�V�9ߚl���xۇ'�n�݆�B�p;�����n�X����j�ߩ@wi�M�����<��Z�����m��%���=ǻq��֩x�):��y#�z�J#��Ft��Dv+g�`)����� ����$�"�(WWV}�0Y?�}b��}�?n�{o�@x(B�0�/nwu�%�h���Dw��
�{%
u���wl~�]r��Z�hy�駉h����Ơ��p׃�{�v������n�GQ�����'�3�j$�#�6�An��p0��3�W&u7T�Gi6B��?�u���R���N�^��ƍ ��j� !~Q�^ZlM�����h�GHUd�ys� �+�^R��=�|:�+�*͹�Z u��,���\�Q�xo�o�>â���ⷤ���춃�U�����������~��}5����\����<�B����q�������c+z�p�8��&iX�4u!@�I/��>�� ��z]�Rߒ���okFI쀶
US�nuYZX-��������[w�y����f�x��������6����e�Gh!-���F=����:_e�3� ����f/ٝė�iU�%��L^6�c;�UXT�����V�ci���S�.]�һ}���mu4{�v�_��v }I�o�AޭB��~q�ڝ#�|�so�}a��v!��7�-�v֕0z��g�e�*�Ĳf�M_�|���}������-olK�����˿|�ҥK���ﳞ���L!�m��}�o���{X�n���WV�+i:���:c#2:�w��DO�����1O#>��Z�3����{n߸)݅�SQ���ˏ���[�����/������?p5ο����W�����9����IV����[?�Xz|�;;b�7�Z���Đ�Y�ٍķ
S�����3�eб��K�1�P.IZ��������?��<��?�{�����G�_|�s��9r��A�{(X:(��e%{M���Ÿ;�3�ό�����4��O���j�<���/34Qsn@��ӷ���?���796N��dF�$�=|�{b���^{mqff���.܏���������	�������'!n�D�?T�B�{���ɏPj`�x��5*����5�J�R�+�&��ŝ/��!Vbϸ\-��s��ۿ���!Ly��իW��g?�Y�s�oz���F9��\�q��?���~���>�~?b� pk�`�G���V�4VI6���]c�Tq���{��w��\6�y?�g\�S�#�<^�ɨ�p��cp�:��Y�_���[Z^`P�"�W^�N:��ĉ��_�:��~�aϡ����^��s�����e�s��{�>�����㫫�������|��w�?/,�=鯷�E�N 铸�%��wÆf�!wfec0����ګ��оë�p§���|Z����V���l�\�~�����-&Yl�����!�G��L///����{���3�����/�۷�ݙ�}����̥i����~������9ޙNg��/^|�W^yȟkr�a���oܸEǲ2���U� c����k�E`I	�}�>�t������'��.���:-���&���ڊ��U�r|~ֆ�硇�P�Q�����H8��������;K�hy䑅�gϭ�Z��u�Cz�m�����{��n���Nz�@x,��y���-A\�F�b��'Et6,�ì����(��U�b����Rl�~�ww'��㓨P�H��aX�It3rCϝ������X�QË�)O�G�g��ܝB���M��W�\IAp8�;�Z8�,�j�F�,LmF��I�(�����s�>!"�{�O������;�������{�sZ t0��������3�@Y�-Ęx���cǎ�($	.�c�H7r��7���-��p�5g�=X$c�	�'3�%ʠ��qC%^�KA?����`��܈q}�(�����ʴ���4���"D.^�N���h���|"���X�+��'¥b��Ik�vx�}Fؔ��+���6W�ǡ��ڽ���. y�6ccВ��v!����؋�������n�`�HTj��؈�8�{�'ǲ���V*�Px*�m�$$R!A��� "I	��+W����ʤ���Ά�67b�K�W�`8�/,j���i�ۭ����G�?ظԉ3`������cAQ��M��=�?�Ҳh-Q�j�pT*'�H�������a���·�?��=���</*P��x�w�{�G.;��i���Ӱr7���
��e��@�R��I3f������P�֣����D]�+��e���1��~Y�h� �K���QEO�K���W_}�-UQ��ȑc��w��o�F.�[��M}���?Gt�����k���G?v��ַ���Jd��a�VC��{��g�`����67FC��k�S���E��kB�m~�V�����]?I�Y�4<�X.��9&$H!&����ǎ�h�[w��Y^t/#�o�W����O��O�'�p_���	�����1�C���;"��1��+����g�Ȋ%Tź^����Q�����ҍ�-<e����i��������6G�i�sE��D�I��0�CuZ�x� ��u)�66�3�j�A�ϋ/��~���V	V_�:��o��
|��̟�ٟ����#��{��^��O/���M��I��V�;.$�y �0~ot��x�b��OV����Ԭ]���^��ZB��d������ģ5��q���k�����a?p+�[vm�A����.��X�kZ�wsFí�0�~�h�mb�0����i�e�;l�q�\ص�k/G��n���~�Q��Ӣ��tiw:O�	B(��w����e��9R�l�����x1��˚�A�:}����?�SZ����w�8=�^���^�"�kb��Y�G�E�s��D0�,���Ahǖ���1|�:����z�� ��Ƶp�q_�a�ݏ�`�g���t�~� c�ȕ� ��˪�$���|~��++�m��8������Qt�6��P[�a�D���Ė"�C�y�g ���{���5nA�[&�G;w�	���|�n  �&��,����8y�$-_s0�H�C��Df���e�B�X��CÚ��pT�{�A��~;���#��SV+(�)����4�|=���m���A��M2\��E��n޼Ξ��^�)�ҐU_�h�Rd>���������;s�4� ��*�v�z$�����=����6����1@� 2pH�p^X��B��� �<�����(8�����5@�x�87���\��@@����?8>��5# �����f����T��y�Y�^/=G�B�e��u&�@C����Y�Ÿ3w�(�H{D���r_��ЯΝ;G'��>�9rp�W��Ur38������������8-�T����b����nq^l
�RPv��2�p� '��W_�Og�z���g�C�7�7���0��
�~���+6T�ݷ�<x0�jU��Pj�O��Wb��
�
�<x��}?�D�L�Xk�V抾��*O@��u��Q�[�t�ޚ��V�]��T.E��k�O��uG�=ąa'�~A6���L�bp�J���=>��fÍ{"^����Olp⫞a�<q,���yqxۋ�c�s�U�W�"x"��+�Y�n�����$n��&����[�v��>pc��r<@�M-`�k�c�?�����99=��+��OЈq�*mh�5[����dZ�'��v�deewq>�� >��.�6���~�~ry&�]�`�~���̈���)Y�ٸ��0���^ � �z�gxp��?��1���r�E������b�02�8�S��q�[�tCp?<���ͷ^��v\̺	3�;�<}�x&��00DWz"�M6Cͬr�	��}���؊0v��j������S�B����+��z�n�]�d�V50o;k굧]�����}˴a��'�HX��>���^mՖf���X|����gB�2p�?��Dr��q�pN=z�=r�a!����;��)w���ƛ�Q�{��gh0 l�m-,���0� ��g��	#�D'��đ�xNLdbc+���8��0[Iv���۟���/gYދ��&���N�מ=�!���݊�\�5�4���}�6�8�.�C�tT�#��[�L�+b�������p<8�K/�D�
���iǸ�@#��k�nG46���������K���u�����N{>{~�7ۀ�Y��hz��v�����EJGG��<������">^�[�y�����~+�z�=LԲ���{O=�$!IX<X���|m8[�k��{^ok��P�
u��m�����BL�K
V �zfE�CB̅öaY{���7Y'��D,�(��u�?��>�_����hٸ����1W�\
ƀ5x1�!Ӥ��S�<�h����\JlR����@��C�wp�6�5��ovhL�Il
?]�#����}��'����5`�a��	'VݵkWiQBla�m[D���l� p�L8��O~�`��j�"�>d�)�J�ī-8�k-��� �_{��{���-�k>K
>����	��m>N��ͽN�����Ë�eqpv���(7��w���{2��`8��kD�gD�6nx����XM�v�����Dl�Sy0~����P�m�a�ӡ���g��C���E�^N�I�� ����+m����o�}���3mHha@dJb1�e0�q\.B�cW�C~C>�?�UN*UT��T���8eG���1B	�� 	�E�ܭ׷s��o��1��0��9ԠY���~���97?0�n]3�
砢ʞJ ��f  AY��"h*}Ybù��� ���e��8z� }o��g ��:��`f�4@��"@��t�k{\MA�m�@�9�{Bz����'~���|7�k��R��z�vdM�����?u�ȣ��	���r�r>1�ʥO�/ryO=�_| @4�� ��>߫���z �I��4�ʩh� +�G�k4�=��C��D�8>"c����A�+)x5��֩<<��W�ov������3K��߅�s@��s|��j�V�������V����+F��DFV<y�#M���Ϯ�R�O�4�F���/eYZF�����F���w�x��O���C$��i�j�È�n��}C��,h ���t9N���d��y�* 4ו+o2Lե=��c�g8&����^��4B:/z�5��r,�^�~'̼�{����������Bc��������*��"E߽A�M�~2�x�A�Ka���L��d��{�sR5�0����p-�����(;�@����b-%%�L.�:�Z��޲ӊ�@�ԣ,�����B�� z��z,�O�B/^g��=|�`��Y\&ua�v��}mņ`7��	����S�K1��0�X[�b����ʔ�UD��T.y��= O�+s�v��k�W�L��x>�hߠ�#��a9ԑ5�]�x�E���^T4��J���ȫ�*�K�Fe�����<W��F�
��J9� _�u,��Pd������?|�`�ӥqR�����xj�g�٬��#?�
��'\���4q���������`X'���U��a3h����.E܉����h�U�QJ�0�T��-�r�I�O�� >����%:3�f���8��������ېW��H�U��,��;=
��q�!l��c��#��X�ٻ��&Aof�������o�ZF{S'�|�V&�D�fC����D���0�f��=̼�*Si�&L��i�I��l�����̜X�Z���y!��n���8(����v5���� {�i?�50�o ���]��z������r˜ '��uZ�ߏ�^*k��C�O�+����l��Ç�>2�I�\�B6�C`r9P��sIv'E�����GH�|�d��Ų�&*�D�z�c��+N>R1�8�NO��l�: ��9���zs�~m�>ͥ*��������}���;bf�tɒ�� `��/z��}�Q5��Na���Z(?,�~������5��8��9��N�Tf���L!7^ߑ�{��#RQT�G*�Ʋ�	�| �(i���;� ���bT�t-�R�T0������A�7fU�~���Um[�����4�5+�����P��\��O*��b��k"L�<Or�p1_�i7ki���ߘ��j9ނ�G���6͸���7F��r t���������ŵ1�z�k�л�Iֿ���jBw��G�c���4>,�:�7P�/T�� �
�t�%K�Ig��t��T��S>L��]�$;�S�<`�+�Ic;|(�H�F�a��k�m3�M�%��<7��TM'pCN�KK�<�|�@>(� ��e�0j��ۨ~]��7&/��5�kTt�IM�
¤{c�Q��}o���y�%;�sr2+
.�J���S�Z{���x��[����M=��pDj�
��9G�М�URh%�F����+-//�Ƙ�j��v{��`D���B��d�w�-L�0����wܲ��hGp	M	���~T���*�E�(se�dF��p3�>%�Rn1j@���h�����N�'�<���f�<y.�=��h�Q�o�l���
R!`��cfW'NC�}W8<]6��T�)�(�C(]^Nt�����4�;��ɇc?��}l��u��c�s�eRj4�*�32�AC���a��Ro*��P]���A��h�5z@�ۙ�O�7T��T�����/� ��|��p}��i��o��z�y�"����HݭcX&� *�熡a~��/���y_][eme6v;�8zp�[��h�y+i��f�t�-�<>�v	tI�2��  q�[䲌�3�
���0�׶9�L�Z�걉�dr�T(��q��Q�$��aҩ�o��z!�[��B�'�s�Q�&դ���r�khOy����X"Ӣ K�%ҚH��d�	��!��ܟ��b6  �dq<�-�t���\��ڔ�H��-���q��<�_����*���p�ٞ-|��9i�X��e���I���>_��C�CO��+�X�Z�Rt)-��6���Ԍ�	�`A#O'�0���)���k?X0��X+BmO���SYɭ��=�F���W���磷`�yL�0� ~�(o����8��	!�)� ��"Of�)*r�:�P\���W�w:�
�M缰�N�l���PE2��n8BR�A	-ɭ��s��T������bӹ�2��N�"`��e�]���8�A�M�ǎ���P��x͕k���+���."z�j�iZI��HQ�����F`��.�����͜I�H�g�z��%�*���<j���I���<�����׃8�k@ � �u���С��n��?ȥ�o��/��A���Q�YMK�:�
(:.����oO��qq�����w�����ƕ��Y�k�ֆ&�s�廬�ͨ�!.�H��:ɻk~N<�أ�ر;�C���7���o<+��](�2�������m�_4�L�X��0����)߰��J������'��~0V{�f��J�Д�R�0�Ȩ�;���܂j*�+���P�Es$����K7���w��h.�"�����$哯�W�h���b����]�C7��}�㳏=.ڤ��s��^�tQ�I��9����rs�ny�5�[���������;x��x�t�T uqߛ�g���8��k\ٰ��z�f�>M�*	VY�V��\o��E��Á���$���pt����&���͌�"��4U�̀I�* ��Ɲ�^:�4b�����{D�z/�}�ŉ�犂�옿��|����,5DIt(��}����m��ffľ�{������~O�N���9���;|;�:�'�y�<���J��G"`)���ĸ@MqBעິnQ�>�дSB؟#�r�Ϸ��^C�.AaƖ H҇9v�����l�O?q�P�ϴ(R=x�݌s xbc]PZ�b������69�qϛ�PLϨFlԣ�T��R��HZ��R�h%�Q��N�Oh&���䣑����T�Nr�j|2 �е�j�E"�ǘ\.c	&!�# B�=��޵kK���뤉����>S���E�i(���!J<Y@��J]���qm���*�MRꞨ.��������j�E�O^mW�A$_�&�͏��L��
���T��@o��k����Uq���~o�SfH�E.0N"��M���Tw�M�F1�Yr� �����ϦR(�J����33K�]A4�4�>k�o��1�7��9�k�!��@_�c�A ��AO��:
4��J.��(��b��_�]���"�a"�w1�F.� �י�>ѐ��#y$��\�ڷ�Y����\�> �&+�q%�vk�1���ծ(h邔q���!=�7<�c����e_���E[UV��[=х4ݞb���;�c�Ǹh����t� >n��Hym�K�W�Eչ}8<Ќ�/¸&�JU�œ�noM�����e���҈��@,鉱S���[a{��%�4x�}�Z
Z�M>i���i�0�U���f~v���F���@=��uf�ut��u-���4-��D��	Xf�hޟU�EI��b�OMuzq:���7z�7|ʊ2;BgcB������ZpD�j@����G,][摳���QϪT� �j
e' ��j��(��Ge��z ,L�ך�M��a(I
�e]Vg�r���t�*�����Զ=�B������`�BF#]�h:h�,���Y#o�󞙞���$fR.T�d��3�[��� m^Y�1�G�G�������q��1�N�-|��:3�ngf����u~:����M�v��HHU�T5��Y����Z�Ҡ�w0+��"�}+5�1g0Н�\ �#����x��-QηN]!��)YB��sD9I�Wc��r�>i����;�@E0�R��Ӎoϴ`���4�9H�9B����K����!'�m�޶t8���u��o9�ʠ	ɷ�� C�����=�\��������̢NR�q�=�Y��&��A������J�ڗ� ��q܈�	���bN��\7pK:��ov��ݍSE�\8q�k7<�j�ͮM���5�T��$]�D��
 �8�����@���;������^��u`��#��`����.|�ї09J��wRѡ�" �:y��:]�Q�z�����rm�
D��[��e>Z8c�~��"%s9�-�{y���;L�ghf6�d��;b��s�NZL�cͫ�+;��.h���/�s��f�f^"�՝�1��u���ɳa��+K˻�;��ϋn������z�����(�c�۹�b+�X����ߴr�葵0�ٻ��oX�A6|��X��0 rH7�m(HF�US����1p~�z��bG/�8q���;�ɋ_����=���3���Cז�2"�#���O5�d���XED>8t��[;w�\��	/\��giei����s����& g�c�G�P��	j0]8WH� �Ej/����ٳ�Փ���ӛ��y��s����ON=|���#�����=hh"���]'U���-	�!
�z�؂���ێ���'��ƓO>�ӝ;�V��N	k���)FtY�8H ��/�Mɡ{a7���n%�3�ݻfE����t�QP�j����*��W��C�<E�%t�S�̱e�,�\Y�Յ�|\���p�{vn8=5u�۽�SSw�����������g����|���l��&�c!�EIJ��DɵcsC���$�n
�VY���o�/���~���ά���|���~������--��&�nt�RgF ��{a���s�^D�J)8Ȓa��R�v�u���W��O��=|���_|mf���{����p�d�<��q�`jz&��$H�Q�!J��x��k;w�Z'��	�Q�3{�����O|���O�Ĳi�#�a�S������=?77����=(�Ji��rpy��W�)���Ȁi'p���ۍ�­��ue߾}t���g6\��?�������O����:�M~[�n��ld������(NAPkO�za��v�m�{��ǿ���}��ѣ��:�|�j}�J��+�y�Ň	z}�����޽+��u����x�37ۧs�:�k�۝��i�+d�S�;���>�g�����=+����z�Tozn���g�<���K%N��Lg����+W��Nv��Y��X����?z�F�d9�Z��욝_;v���ɓ'���l����/-�:u��i��Ku�8�Xy�� "�f��
i��#�@�H�}6}[j������8����]��:��N�E�q��|�O��;�k�+�?��_����f� m��u�rW�㎥#G��M�c����n������y�嗿�y��iq���W�����˗/1J�}��<a���w?s�'>��!8Eh�tZ��w?�f]���ѓ�.��替&�~�̹y�]�A��_��+W���q�~hK҆�w�q������j�T2�-&�p<����}_y�ᇯũ�ӧ;�!��)�^7��K��ݺ��ս�fs�̚K����ǎ}�ɧ�|��W) L��=����o�R��-�e�y��ϒ���Ad�պv����������>�f��op��z����� X\B_�W+�gf��p,�	�Mg�|�bY�↯V���s���l�q-Ǳ����μ23��ÇG����׾�wLF��УԶ,y�A���߇�=��Ӓ�b��C��+</�^�	 �|���|�%n��di�S��{��H�"�n`�����̦�a��L�q�J ��y��b�
aˢ�Hs#A�{��I�l0pS�����#���IS��� �����l�c:Sa���A��cڮ�S\����v4Ѿ�	�-�4��h��ܽFZĢx���Z�4�����\��)��v;o�Zc�\-R��J���f!�c��˖_���ZS�4N%� �9L��q�GZ��2����E��� A����&��e��yNT��8��P�r�s�A��,m`��)�T��c�h������S��c4���[�ϊ�^-����F0�|(�MH����m�|�!v��]������{����c�@�s#Ij�`}QN�׫�'k6�8��6yI����� [|���i�I(fCN@��/q�A��Q��@b\�g��Vӌ�)�k�}b�@i3eˁ/M�</dY%���Tc;�q��i�pUP����H��#���������+�(�`.�P��7(�H�L� o��a�S���vvp�
�54m9dieˁ�O�{�e:5
BZB3��=6�|	���v�+ ���"��Uu�0�F�}�I�bȍ��2� 
Q� ��y�nv�٭|l��������~T����=#X��f|�qD�Ѯ��_����Q��# �:~X�{�6�#��tT�LU7xS>v��aw�n0*��dY^K�>�^�����&���r���+,�f��a�h:
�:*�J�E�Y���~��+X� ��'�kԍ��{�}�([|�'3����a�Y�]���c�
�K{(�(�/��Z�H۠� �$}��	�M���$���&
�/9o�u������m����n>%z[Z��U����l9�!p�+���\2a���\�k�+�|���*�_�$���|��x,�%�'�<�bjj�h��I���9rdl�H��DG^�e��H�W��Aq5�,&�߃l9���/n(j�N�bCۖ����J1����
�B���ٛ��Y�EL�L��߈���)���_ǉ������.�AH~YT��v�����||lz�$��->��B���d^x�n�Щ��D��#�T�e�dwk���ІzS'�) ��$	4�m@�A{ Y�(��D���5*����,�jI`�_�����4�
C�����������>h$$y�@��y��ؾ�+��r�͔�Z\�5&�嘪��\��%w!j��&�P�r����e��a�-*Uɑdl����AcEG�`0�=�W�p�>E�.3�7F[M��mv'E��T�������1�����'�=���'m߿�F������w���&L,۱y����n��bXCJ$q�:�U���k+=��
�����@G|��h���->�a <�Yg2��֧8��Y�r��>;�%Ϸs�NI��4z�j�fn��ʖ_�K[G�fxxQ�U �D�dn����H�Z��'@�W"g�2��	�->ŹV��t�-��������Q�y�4�hN��XOC��s�(*[|�v��jj/�����B�;��v�ˬ�3��;�I�a>�4v�y���j�iU�?�%��=�L ��WvsD긹��������f̔�pG��[;a@&R-xXtϮE,oG��"�%%i�������)�a��uj[�ni�������cȉ'���G1:�4�Z0@ %&T���(vz�����n����j�Y��6v߮�D���S�T�l��/��K	|���͇}ۚoRM7I�G��\KX.��f��x�7R���B�v�,�CQ��"|��_ͪ��S*[|�F���/q�����[c�/�N��4-䱱r���N��H��U��� o>�`c��N��^�� bD����N^[�$��-�~�����$�|�r- �����ouԢ?4m�oR�+dj���!�w����,N����$�h)��8�jDj]e0=*C��Ռ>�v1����״����A4��~a0�	��HB�r����S�Fl�����6R�_4�`{V�$�@�,����*riI���H�������ƫ���Z�Pץ���A(AJ���Ʊ�����H��6E��&dZҖ��]8��s=#qy�*���R��)��=/�q�	E1��$�N�L�h^�����ة���i 	E�Ֆ �\e�����"j
=�YlI�pcok�I�I9U��� �.t(��j��� &Ǳ�ly8��a]�<wA���D�':��l��21��,��k�D�0�0��r�cK�|�� ����Y��CQ����	כX�ǲ����.�"g��h�gv��	 ����:���\/A�E/Ŧ7O,�t��O-��y�Q��Zn��ya���E�ܜ^XuM- 	��m��D
7Ș[�&&T��B����^@Q�F�q%d�b�
��ډ�QQ��橃c7M:}�gK�	�->E����n��dՒ���D�42SQ�G�n]+�>zfP� ��mב���d	 �0�th&s=��ˉɏD�74�l���I��#��(���*4�#��ߤH�eҵ����]��d�6�خ��@ 7�u�|���?7�d� ��a�[4��̓"䓡�u�)��mٹm岮!�t@�x��b�\��<_���m�k�������Ońʖ_F7+�2"�)F�/˱���z�����8�di�v�]��ҧ ���<=��ݻ�7++�G�س��W�hX�Y��eˁ϶��oLOO_m6�A�|���ql������o�SS�v{�\�z�Gַ�cCz�3˽^����.,/�}lee�;?ӊ�P�r����z��[~x�С��ј�8���]�8������/������o�o�w�~r��3��q|t��?^^\_�^�zu���'߾&&T��N�<�����v�n\!C&�`=ٵ�Z�ٿ��e��Vw�Z|��v�[fW^ j}����fɖ �>4��5�ă�Ö���]���n�    IEND�B`�PK   G��Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   G��X����H   C   /   images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngC �߉PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK   G��X?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   G��X��) oj /   images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngĻg\S��=�2�
��>zSzG�w�BT���	�����N@z��	��^H'z �����|_�{�?~��疳�.k�}�1TS]��������\IQ���z"�k����Hg����\I�O��ߟo?���I�Е���������:�� ����������ks"OOOk[W��N�<�.��(	Z"���d��x�m�{������O��݇D]kg`%��1�hU�O\dq5�Zl��|�M��l?���c�0*M���Z�ZwN��a��j�ߕ��b���������ad�~���ޒL���~0,�Ƈ�/�7d�|��b)���_N�;��3H�xg���c�AA⿏eri:��>GB��},��i;�w���J����S��E��ٮ����G#�%�ܨ�1T�{���''=���']|޹U��]�b�E�џ?*�������W 
�_@�O㩤0͌����g��A)Z,��m��ąO�s��V��I�k9y&�+����u���58����|������U�J�t�ر�����M��/���;T�1yD2���k�K�%�$Uf�U3�W$��B����K��"T?ϗTa�:�
m�p<k$��W�����YeZ��<[
�7.�����5.����/���y�_���L�܃A����d+�̿��!s��!s
�W�B.�@�r;Ku�&bt�����4��E�Y)!S�!��,�c�����aAX�J����e��[5y���F�,����f�i��x�d!H��y7��<�_�Mv�N�Q椽�Ѹ^y��-9f�q�~�q$�W�
^5?�]�?C��5(��`I�VZ��4[7��|���H��[��S�M�_�ߞ�x"+P�
*w�M�n,5�p�?��}���y{�|y��omj��M�z���4ŉu[_��'u��}�f��!f=�J/��do���{�+��鄩A��bKw��|�1e�&V�~��I<G��t�1[ˉ)$���]w�ޝ�.Γ�Y�"pi�s���O��S���ſ�2�Ϳ6��]�F����n4JF�y0lM�C��!�ު�(�AX�o�֮�Ue3#y����ٓ��2<�`�;�C2�Q��J ����N��c�u^��a�&I�^7 BN��pJ�G��i���q��	�j�tǉ�z*�?v�_� 5�[���W/���)��6mwƌ��%-[���8�.��'7r���xћ!'6^�h �����g��NS��%gvu�sώ��.��7'$���J�L��}�S�/�}ٞf��|�kb�W�)��ء杜�>v�zQ{P�uoQ=�����d�ꃀ��b����uM���պ�X*���`g���s���㍋�G�G]��H +K��,�	��RC�T(��3;��Wτf1j��D�!�%4[l�w&�e+�:��zI�^5x�2y�A�9���7N��e����-i�w���[���P�Ն'lE��)$�ɏ���S��0�a�!m�� �`D1�װ(\o�xoz力�׋��D�߁ԫ]tg�g؜!��C���t6j٤��� ���Z�=_���c#�_Q3��}C ��$����mD�$~�-��I����8 ��Y��3( �s���6q�\�1m�Rc�B���Wu4~��Ū��h��2��z�(|+�q���9�h޷�+9[]�TS�vW��e�Jr@rB�g���/[a�W�1Z��������DeL���O�OyD��u�ԁ%2�(�����{�F��lk��L6M]��8�z��T�B3�x����Ⴑ���gs׉ߙ-�^�6/�r�O�CV�3Z)�]s�P�!:�۟����C��9j��Pa�2��l��j�b���Ml�	��'9E�v7>�o��V�1���u*!�h��ίޕ��	2_G����v����X����D^��l�I�YH����z�����Yr�I����g�}Ӫ�a ��c�Nb�wO�ݝ?j<������Ĵ�ZN�]`�
(��3�i%_�F�s�� H�U\�fz��kw6��w���fË��9}��X�Rx��e�y�d'-�� ��!��;��JL}+�����S�{9<���a�0%��i��U%/�X%��T#��'���䡚��3V�[��)\f�3�H�y�Y<�c��j%��o���vR��F�4�=��K����,�ұ��؃��`�Dim�i��b��nNT�d|@yLV&T�-<��|�K�1��#�����;�W�s�^���]p�髀K�ـO��.���?��� C����kLLH�#N�g��oE��NF���|�e�����!����	�W1E�!G�%�^=;Z�f-2f
�36��.{6N�}�S�;��V�#�A��އ�E7Hx�"t�t�m?<_՟�?��D2AkMb����P�Odv�.r���c�"�x/��|m��A���f�8qr*�����b�u�����W3%^L��[8�Y!Z³kG�7k~ز
�:�S�)
�����l�c\A}�����L�׵�o�Ε��`,���|/��K�G]צ��h�����g���s�f,��4��e2r��Z~�>�Do��6�C|v�g�u뛳��tb�CeOw��]�c���/i�t�L�N��{�7+?�pя�Y�o �W�g���u����&
F�fLd��o^����>�_>�����Ċ�/��Y9dg41���w���:J�B�s��XG��+`�<�vp� �Ê��2�&����!,��nw�P���ك�-�|���n3�{�����w��|:�n�Ȟ��i�~ʑ���;�l�}6)R۹=z��EH4�_��W��'�5���.��A컬�l��_�p�}�����'����ض�Lz�VΥ�/����ƌ���+��J`�hZN¥'ŐS�f�M�ӱMz]Ig�Y�8f��]9M�Ư`�SR�`l���pA����\����u���M��#g�!H���Sy��fm������CO�-�����y��U�&��+@e�Ǐ"R�1�4��T{{����LZ��Z�ж/��}���#U���m����:՞��g��ɫT��k&N�詝O�#z��"{!�زw2�n�r��<8�c�]jǼU6�r��r�>�J@n�W*�U,��|�i	a����˼��oB��~|I�X6�h*k:���݆�Q�G�M��P4d�3s[p�Uk���qc���X��ں���cCs�J�x�-R��tojg:wt��f|�9=�c�a��s��J~�RWs���E{"U�G�����t��tj�*��
��1ũ)��1M���ԫ.=��T�㙫�
����q���H�-u�H�0=¹@ؿW�Y1��JK�:�"��J�\=LJ*',=�g�G_{���I�~l�b��w��G�\��Vk��=�juڡq~�˪��:w�q.��&*XUz�"�Ķ����ι~}kI
�w�2�^��>5u��?5}��%N�*�@R��}1x ���4C+�c�����i�Խ��*/��3����O/܆�7�[_��W�).~b���������72�}_0������-Zluq(���*�Cb(!���G��.8[�~��ɑ'�y�#�N)Sh0��wЦ>��� 9�` 4%�	�m8+������� ��W(��Mlg��f�z��D*�-�ӗ������>t�5t�IO�]�v_w��DA74K��u���^m�1��q�6��xp�'q=%����AP^ݘ�ݸ�nt�t���t7e�Y����^r�]n�b�f��[�¡9�o
����8^հć#n�w4��*�}n(���r���Q��U���i�����8}k㟜o�ש�>y��,�;Ѧ��b�y��]z)�����Zo��n[g4�zٚ��ܖ��i.��[8��L��1�r
&p��{��2���/���k��G�I��%0R�ۘ]� f
�}jY����9�a%�2��]�0�Q�������k|�L��&�Txlʹ>��t�&[Y�ar�}˰�����F��q���L&������;���/WdГ��Z&��N��|�d(j��-b�r�^Cֳ����ܖq��V���|҉u�:>Hf*��e��벤�YZ�3BS�����|JQ��!�6;^G�#�g	>�v����L��yºL_�,N&"�����u�Q����V@�w! �������m�*1�S*,N1�g36�B��J�=2�o����/�
��L��}H�����\��+���������"NwC���-@*�+a���&�({� �����x\!���ԖJfc�ݧ"lL�J�R4ob�.��}���I�d���d{�DB\�l[A.�k�@����0� u�D�	��y�	��	w��[��^'�r���	�ƎިC���Y��B������/���P|��t��y�d��Y���)^6�{�:v@��t$��|�-�&.r��>� �L�zGjv}�	���OgFq��?6jF���)�
��::ߝ�^*���Fz��nOn^�8��W.ǭԂ��0L�:Q�7�<�~���7���t���эh�I��?�@E�?�o���v(:�����5���󼳈UW��P��Ʃ�8��~��h��YN�r�Mi��BNW\D�m}�θ��a�c���������}�)z�l�j���-��1S�;ǣ���л-�`"���$�.�x)xi׵!�rf�:ޗ�vhVLdc2# ������qiݵn��C����7"s�#�Y������lR�+�0)�Cݷj�yK��I���TgҮ�䮇'�a�׭=Z��ўL;⸕*�����@�ƛ�~���-�-&JL�ĺ1�bC�D�r�0�%��~�g\�3���=0�o���=}JEE�ǃ�3����'�/�p""mO�6K��((;;���ar�瓼�B�r���^k�����7���?�\&FIg	|�958*��Jζ̩�GV��!��8�v7�i�P��jɯ��z��p��7}/E�A�W�y����ѭ��D8e�S���1�]t�|v��w�v.`/�Un��;�U�P����2�d�����;tH\R�4l-=l��dZ��(��{��^�-��2��(���0��0��CF���������J�--���޷�_h�M��I�ޭ���y\ ��p�*a�;z�K�G���?S�B@&r��RC˟���v�Z�$�\v^��I�܈n�;[��W'n�~�@7�> �b��4�Kdq��[�2|t����蹃^��6�JRp��@XES#���?G��:�{�*/le�W����yI�u�	�~���VXכ��
����~Үk���['���1_3kO(h��4�Wۍ�$�ac�|�>e�  Ks�����'�c�6w$_p�1���c(�����~Y�u~��i)lG��k��&w��',���B#�ё������m�u��D�!)�]� �>�Z�2�>�fM��-���d+���v�����+��(��S6�X�B����"zLycC�рLm����7�U��0_��l���~hH3��N��JD��1aP���}[z�W�^x�Rt�;��<g��2kS�V�g���W�yꞶ4v�;�\'��w?e�۱�]C��{S���17�Q�L�����	�Ļ�y��\I�y7F�)�uk����X�D7׀K��
�yQ
��ρ��rXpm[[����$|<{�ߟ��:�S- ������� Pe�'|�uF�*:�"�6��h��6��w����:��=1m�ß����-��"7AՕ���Q��/��s���ve+�/JԣM`|��f'��@����� -��͎̀����!�w���'�$�>@:= ����F�Syy�3��D�\	���C�ʒ3�� ?_�U#���g]�L�2��n�~+}��ח8_�o��a*�X5nSD�w��s���g�"��~�i��ްO�mLs���l��}�WyV=�^���(�*��c�Yy� g��'l�Cl�M��X>�U�.�\C��+B���hi	��v����{:&&�[ȭ8UsC�@�L)�P�6VV�<��Bm��y��JߑXXі�`x^Ͳ�Ӑ�~���x5Ke�޳;�F�	"��k�BGJ�,�\� ]���b.�aC�ً.��s�0��r{_��8[� P\ķ���������ʠ��+���f��k�a�ݦ��!Q�⏐
�pAMދr��k�&��%3J�7~�%��f�n���ښ��.HI�U�@`3�[���޷~���9Z������{=��۾�i�9�s����k=<�7���8����;�!�~����\g �D�筕����~^ѧ��{��"�H)l��h��O4~|�n��?��d��a��HU]�A���L�k[�]���_g5&�V�q_�|��S>g뭿��a����U�����9
���vp={��O7���u�ѯrarّ��ѓ��2[%Zmk��_O�l6-2YTD�f�W����g�+�q�w5�~8���8�nD]�V�Gv�3"9�,�M1ar}��m��E����"�{Y���Q����6�U��U�,ܒ�#���t\�dU7�`f��ҫŴ����0Om�e�:77��OC����$W��=����x��{ �X[~�2�f%�8xO�X�[��-ADV9o��D��%#�G�\�3�LR\V�c�N��}������Ís�RuY�\;2Tb�ǚ)��3��V���I��
Q��'���5���F�&
��$'8�f���A��ɄD�ۑs�I'��𻛺ƵVJ�M�?��U��Ǜ'�1Hp�<�Rݠ�U=b_d���)�Rf_�L%|�`�=�]���,�+��G��&��F;5�,�Z�I_X+q�Ln��ޙ�~�|����vT�5�S���v:�P@皂�V�>ݞI,Iٔ�"��%塡ɬXNgh5�w:]ۢ��A��*�*����Z@����H�L�;Jt� ;[ ��4m���N��6y�U���kq���7��������8��3�m?l��'ޞ���j4���g���b��s�U���97�|���`�{���2�1��]L���)�6��k,��Ї�:å�ۂ�<U\*�55F@�3Y�_\T�g DD�a���ɋ�����\^N�.	���^0�^�R�����L�c��9��S��I��}R��ӭ����iX+���~�n��˵�
�/c5pgS�r���9���e2��!�=�#��W��j������r�]|��>Y7�\V����ɪ����[��m�J����u� �r��@�1�6�1�ĦX�<��`�e,2!~d���ex�b��`�ܨu.�{�h	�2�9NN?�'�S^B���wGa���3�9��ɺ��PBo�9�ae�Z�^8�(�``��e� m央�Q�G�T�a��� ܌���Gg]0���^!���k�+�U>�kvWx���l)��&�X>��j��7��e&�<aw L������>��!���S��B�m��G��>!]��ʟ�j�o/�PQxQC
e�/`jS	?;l,07P�5��a�ѽ4���o��#P��bwȂ?[�l�q7P��'H��G@���_nشS�FR�ZJ�[v�vO��q:@��u4��8�3�4�z�f�����\[S��\YCW���0T4z�-�U��J.G�m`
m<����e~LoN4 1�����5��j�pj��#j��x9w�C#SA�����
K-�xN�.�K�i4�o��(��D��٣���K �dP��Ј��{6��@���lʞË�7K��*����@������'������:�*�mp��^���L���Td���
�u� �n{�f�j��)�;�d�4��Ƚ��6MQ4�
AO �|��\ݸ����lD��ig���o���Tk�&�S�q�ǌa_�p��Õ�\����d��aR$�buچ��]q	,ݏ��4�6�5އ555��&`�@��8>�.� ��>�N鮸i���Y2�iP����c��<���p�l��;��&Ӗ��=�	�EB�C+no��Y�ۓ�<����J���*�l��_P�P$j2&Vr62C�ѱ�m�Ĵ�d�ׯmn�~��Ͼd�Y��I�w���H����ۃ�z	ey
�xYH�5AIM�<\�J�Bi�9����SO2���J���u(���U�fC����4�]V�o��������J\xL��j���o��wg���G���tL%A�X
 ��f�-�]E%wa��lq��9�ҿ[���c�]�� 8���I(5��b}c�4����/;8덧�G�џj �~+�6��?�ߜ�,]8�Ձ������U�MTd��;F �$v/?��&t�z\�2@`q�|�?�g�.����Ϸ�Y���j&�%����yԣ�j����F�Zw��C�������c�-[
+�B�aUE�S�<~j!m¦�Wb���j�уy�K�vΎQB�_2���H�`�|mh�:�^���zA�Զ���f��Q4������|���<Wj�o#���zNm&��	ͭۻ�k�����o�x�=��N�pz:9�9Jh5�=����&H��z\�����X��1��������s�S�rkF�	K4?��c����]ߜ��˝��v\���ޙ7s�\���#
I��SSu/�7V37�f��ǣ	���	�U,|'Y��8kd?W����������+ ��6"�]o:<�]�6E���+류�I�q@h���Y���{(U-�ʤ�ؗ�.��R�C��q�s�e���"�xr��/�<X��.VΞ�6�����|����%�\
Ҿ	� ��O�����Te�X��9��%��x��녔n�i[�)���El��4�����[��u��ae
�SVSX9��<�Ǉ��,��	{n48$��K�T�G.�D{{�k�����k�mG;��F��|��2i�m��r!��N��2����.��?-�a�C�s�,�d9��y���G�r��6ڼ�>:w�:�	`��H�Y����l��#��zxdZn�Ď�y��X�:/��&���%��0��<X����RW����s�yK���L[Q��/�ϛ4�6�-_�4W��蓡B�>�ΰ��۬��O�QI7v��fKh$�be�����ٺp��z�����WA�)�����vH�h'������2�bz8�F�Y\
���wv�j+ʗ��LM��K�<d��l	�j��ى��C���&�W52�"�J"B�'�*-(��tR�����р�L���5�"�~�'UjZ��j1|9o��dT�T� F���P��`���.��e^O��Lk���w^;�>�*�=�b�����+Qn�N����Z����&#_��oV/��۩���νKZWrB�A ���w�b��I8{=I2�Bh�MM+��vu���8A�ˉ{�δƓ��!I��풴| e��U�{��Z�£+��@��o��B< ���H���K�s+��R/pn�@�-��cִ��\W:�W�x����=��e�1�g��Y1~���e�$'=~����L|�d�|�~�/����/��̘V[�kmCKe���r}s��_ӥi���+�م�Z2H����v�ϒf���g���b�V��0���H���ݠ�H`R�`9���ۏM�o�z���,U��%G\Jt[�:�Ӧѣ�e5�0�{�Oj����7OJw�u��8}D�X��(?�d&���{���`.ğ>�;��Q}�f3ͣ���&.)��#����+5.�J�A=�o��o&��,V���Uߘ��5*5i�`%��v��z�;Y���C�Nf�D��{�SV9w.u�������ĝ�����f>B���^��c�����!�n���O�*��%8�UO�������S�'��6H�,uO��rG��.]�t*����a�_8����ky��j�琎�
��7�\���/����_*� �o\ҥϊ�s���xr���!U���0��������,�`�.(���A8��H��B��*<����]2v���f�R���t����*�
wqO�F\H_��I��R�;W&�g�	Cq�,|���U&�f�=�"�݁��W13(�����=����!*�z�h�I����Cac�Ϋ�m�C��3	�Y{��@]���u���������LWZ���p��Yc��;��|@l����*�/�*VC�v��[��)Z�`�ӝ]��y���׏�ofl��e5��d)����PJ2���󰜙0���Y�Mݳ0��YQ���㟀�^b���|j888X�ZJ��&s���x�P��b!f&w��a�`��	v���}��](�q��<Sx��t�-��
��*�QU˲�]��ˊ����W@��dq�]ۇ�������N��T��ap����4a{$#��ʵ��#�XP�<$���#\@�8�-o=eT
���Ĳ�C��FNx+�+֓}�)&�M��/���8�ш+�X�����!$j�=��{�G^�_ NN�~{5���R| Zvg��	��Q�3�h.X=Lf���ߌ����lQ�=��O��ٚ�/o=���ӳY��,	�g���s���3�M;S3�*�9bS�i�>�OH����3S�Q��R%�vdw�1PX�.����oD�D���a�,�g��l��U��IF����5 ��}N�!�R�V��Չ%��c�$Se���Xy��i�}B颋m.��� d�2U�m���#�)s%�}���ˏ�O=�u~�z����=�81�$�1F�P̳267�3Se��1�,����0��'����䖅����D|�(�l�?�f6�1�����>(p�.����1E$G�<A���p$���t�����w���QNr�nAY��s�I�Q�)A���������F��i��q�H�\+�wi%9n�'qU��%_:�d鍋;W�c�?�q�5Y����k���c	۷����t5ޜ�s ����H��bH���Ÿ�.���Ƈ2�x=��zV$!�{C�r�y�� \��<��{c�_dT���	°�ժ;�py��顺��.)��םO��b̊�V�Yn�Z��0Wre#b$N�k6-�+3��?��%�*��d�!8UH]�w���z�ґ�Q�L�a��$�T�A}����E�\ �Xx����?C؁����bM@:�}����͚<�/����`d,W��(��^:�s�	i�V7�1e�\�c�l��G�
�˰𓾰&��{Ҁ�q����^�48}:���j�=���X���3�ڴ޳����:l[���w�o-]�����i�-T7f�{�t��~�M@g�L���ä������+���(�u�fվ��2[^օ���{d�Y"�0����I����!(��P���|�IҠ	���R���o�~�Q��,�4~a�c5
R$�;�{������Mռ�u�����Z5G�xE�������a�/�?W�UIy�#����@]Vb�����B�OK� �/�����6�ɺ��<x�d�@ �Q��k
�Nv.��6�Ȇ�r��t�۽؆��u�*6�YU�_fk��������C����Q+����6�ɾH��6=��Ǿ���'3rvWk��x��O�.���{,��{�G%��C{.���VF����{� :��_ʨ�J�#oPo0���[��HY\��i|(d��+��8��D'�PKk�Gٍ�jl0����2�ڱ���a�C��Z�km���&�}Z�?��v2�>���߼
~��5��g�;�#P��M	+�1���9��z$?"����΃�M��/��4�{�*.�Ѐ�����>�S���W��I�wy�r���y�^�M�K2 �NP�q��!�Th��͟X);��ʗ�H�`�<ᐾ�[�i��'f^�#�R}z�(���/kE��)7��$��ׅ<��[)�
�֍CJ֖��'��5�3�j�lPs��K��V��aO���l��YO�|��O|r�5Ua; �H�-z�a&�W�sH1�	+�#&~A)�m+�vD�%�U}��z�mN�u)�z}�l��
K=o��_�_�?�OX|��ǋ�`��ir��$�c�]���_����k#��h'���	�eS�e���nB���4�&#1Vۍ˶��I��p��ں4GIC�kc���C��c��8'��b���`k���������F���.!��N�vM�r��v�\>�Ą�7��M���w�Y�f��v}��Sb�'V���͒xp�!�2xUU����a�~V����gxX�.5�S�?����r�5~)��֪%�]{�+鼘�7Ӽ?�Z����G)iTOb������������(.Y��ŋ���P��dڬ�n��{-�	cݜ3��Z��3�:r��S��G��2#W��
��jk9nF�Qc9��lR�]�����[{Ψ�z�?���]4|p2��`EMbI5�B�+7u��fɝWР&'iֳ�7���bl�����<L�E\#h^=��B�����_��;���^Y�)`��6d����֕^����r-*�j�)��p����ϔfH}=uH-����2Ϲ�$&�Y�x}��\j�F�c?ơw�qP��nq��/���P�fs]��.����ݞ�q῁Qӿ�;'�&t���o��y���6���|��X�p�1C�އ�K���9mK�����P=���}_/�� �u(�8/ƼmNV���t�D��d�ed2M�k�0���O�N�)�ք� �ɫ�k���Q���M���js	�vU��7��b��4Ԟ���#
�Gt�B]��o�0OOx���M{_�3tw_��w�`�>v��/w�it���J�N?�2���	�Zi|�:FR�����7`Z`��?���*�Zn��F��~a����{8�X����=]��#zh>�����Ԋ���b�Yj�#�����g
.�RQkB?.����|���]p�g<�����֓�׬_	T������2b!C�E���x	�^�U��/���m�j22gՕE�����]�B?�B%��J�$�j�����,�`���}�4����<ӎ�Z���&O�k*TՈI�] ��Ӟֵ�/XA�=�[�`VN��f�"<���S���ه��b�w��`2��.�X�7�Rm�V͑�Qn����V��x�G�������o����z���|��I�?�(�ܙ��¯t��OΟ/h�ǻmZ�.���j���?���*�%�ʟ�4L�.#���RVE�s)77Y�s9����? �io���X��%�-���x;q�p�ˣA�ҋ��v)?
)᧻����Z6V0��\��;k�( �x* ;NvT��_?=��^3�xЋ�*
 (��(��m0��V�1���)�G�;�Տ<���t��'�m�����a]�|�hq^�N�	8%���Q��Ur�SF�=J1�p���H�0��m���o[5sg[�0������_���^�뽿�_RV��u��	?D��U\���_i���N�0�v3�o� ��~�ɼ�
AR�;�]�n��?���
S�N�\�
�vt.P���+K��?�_�xnb��,ȹ���b�;y��f�����Uǀ7��.���(����HQ����ôh#>b��u]L��a�/��fx��"��L��<��i�!N�e���X��2>� ��V:��3v��QB<���������A��z����!!o�X�\��_hPIE��Ѐ0��}��Gf^}��%��~�W}D�v��t����#vy�Rh�?_e�*�Uv�8Πƞⵝ&1S�6��D���n�$��F2�׳�Gقz:q9��k�3�:�}9Φ��>fmL�M@�V8̏_*U���?�;�nK^��y�-֤�-�:	h>,�w�K�Z ���}iwǡ4Q
u�K���%�"j&��t��O
�6�����v=�8���]\S�HŔ��[xzڂ��[ג�H�$?�Hz+��$����÷�}yt���WC����ؾf�^E�+��Ÿ�j��d���i�]�I/j:>�H�����3�B�a?���ۇ/z�k�:M����N}'���6�<�M{�H���x���.;B/�r"��l������O�c�/�H5OqzJ;�|�bSN��#��0ʺ����z}3�6Y��y���\��:�L�Ld�O__j\W����"WWwwrt�"��3�B�����_V���bV�Rb�Ѽ����)����az,[]`���s�}��$>~E�R�=��=3�޴���/~V��e�g�F>��]��'�MM���Y�|����^ѧ�Yeoʸ:iA}l�OO���~�uB�9_�ڊ
�r����I����ݐ�<��'�w�n��?���=�}�U���EH�%^�D�4-L��NS�%�Dg�T~��6���b��rl�ê1]����R�5/G�#�O���B��vy/��K���ϓ�|+���S65m�!�37�S���S�,�3z�
4p�Q�]��!�o���1��-n�IW)�g��'�|���'������{<��W�U'���K�1���k���kc By���� ���KW��ge[ճW����=�WQ�e�M����Ǽ'�Q��S�����mUe���@�+��ѭл俆�㲲�߸qC�g�q�h��o�ݏ�%��Q}.�T{�
�6�R��|�yk#1#����c�W����.f���Qr~�����}w;�n��\$���=�*��`�2���C�-��x�:)OjiTd�"�>,�}�_H�����p��|�������~V8o�6�^�u��ߵ9�~�
m�=�Xn�Pm��q2xp��h�霺�t�-��}_�}<;"�W��$�bl�q��-�E�dcs�rb`\�󮔺����8���^B�f�.�Ul�,�>�����{���\�ԛ���U�%=Î�`w�zGH��=����8\�2�?cgz�Nã�tx���_i(��ݩ��g�S�� �τ�+�;���P�	n]�ҧ_��6N�9a)!�mu���k��{ɾQK���ڗȑ��DP���#��I�^��b���T�{�Q��[ʥΟK�d��	�h�?���5T{,L	�N�GG~�brS�\��w�xyҼ�_�����F�u��4~�	W�A>�����R)�_ZM|Y���x��D��4��C���N�>�S�ӛ���.���wo'�<[��|֥]��ǁ���<M=�[)�ܙ��.4`L|�N���U��-�Z�Bҹ:{�TGa|�e��������vά�])�:]r�p��3.3�3u=>� ��{_,0����&fͻ˞��&%�/�����!��������D��o��a���)���q���j4����	���l�u�$fZ�_�+���eRW�|�������0�����sc	��Gb&g�q��3�t�򛿼�Wi�7�E�b��$��;���r�U�b��{�*Skrپ\�m��i�u�.'>�0�b	����',>�0�E6�|W���6�P��#�[�%4�O����yX�����2>k�D�<�����uўs�
?�.��-�����t>x�h��rҴ��a�f�)HY�o���;�
ϑx"U�^Ys�H�;�-����C�<Ðk�B\VKF�Ya�]j�u��t+��H1|��i�<v$�]4��S��U�P�9WH�?sn������5�_����bO��~�n�r��jF?�_p�`ۈ0i,w���`[%�����������r�vڤ��y7F.�Ky�N?��c;�^��D����<�� �k�t��}gZ|
���vv�8����߅"���N�_�^��b4j.42��c7h��CL5��K;�ɣ8�w?�u;btK}*��O)\цBu�c��cz�o*N\�ku�������3��F4�?)���ԇM�f�D��O润��')>ʴ�x{5���뫍W�4��nL?�tq��#�6�i�xy���49�}pP��^�+f?]#u\���s��a�1R��'����x�~ay",�e��g̶�'���;[�S��{Mo�ɀ�df'���C�\ӆ}J7�����Ơ){��[߲l)4�s��'��)��UA��ύ@��JAb
����b�
2�ѓ����q�:oi^��y%���q�V���3�Xv�n�^��_��-�1�!���͸��^�P���e��V����n)(�r��w�k]|t�mdP��>/X74B[;ܾ���	@� z�z.Df�}݁Q���n��IA�Lg;�����0܀�9�w�W�X��%#jv������C�aS\�f�������hi(ɯ�Q�5��6$)4�|~��su}r����Z���<r������י-g��F��_B;v20�ߚlK��E
>.�wS��?}�,� :0Z�}4�� �\��)>�o������q�㤥U���<�fX��¨�K��[r��S꘥�ƶ+-��1:�s}����h�(>����1��P'��wa�s�����q-�JӍ��uy�t8���$HX��x�P�o�7�k�U*��t)5�o=�#���Uǘ{������^dOB`n�����3\�� �ڶ�uZ�v������9���c���w��Mn�
�J͸����]܆
��^��7��L���]�f���n���C�[��
���!K�����C�y�|]|�������ѩ�z�5�.�ů5]̆w�)��[�xa��&i�[=����vW��[�ǔ)�{�LX�������\��M{�_�=�sx����F����5��!��]�ݤ�>S~�K^��u3r69��5ɫ6�E=����mv�[r��V+#1_#7�����J�1�,�UFD�ȳ8�ͨgs���=&&�}|�9�w;�Ь�ƽ�A��hR�K-�n���E����,���Em��e͘O�>P����{�Ze��?���q�<���(���f�q0�KV��Q2�����]1'3��K24������$�*6�c"V��\�SέkG�-wwhQӒ�����xX4�,��V���Ӎ��Am^��D���_yVj����}��O[,��1%�@q��Ɩ�Aa��Q_�����y�;~�_,
/�(8�|@`7L��PW��@��;&w��^t#���,��<(��h(G?4y
�7����Lb�I��S�7��(�_+Z���F�0\�ch���z�xc�=���k�$���k�����&�A�CB���A������S	��;�����Y�ߢ���;���0�����\׉*�ݒ��ް⛹6gv���5D�bO�!OҜB�߯�ԐT�B�\߽�l�ȢW�[�Q8���Zk].�p� ���\"�G|Q>~��s���C���Ć.�tD��;����.t����\|������d%N2��4����WxG��]�7B�_���4~���ax���!��BZF�}U#����wϊ7ڊ��s��wM��[NԵ(ԤiT_��4�$���Cr;����b�W�������B���?m�/�{��'Pܕ6��~e�H��{�۟_��L�Gpۂ�Z[��z�YD µz�hT㲷]���b�v�Ma�T�M�9���C��C�@��c��J�KY��yH��x��-�h�\����˒��m�8�r&����~�ގ�j�G�*�d�qB��'^޺�M�X�y�f�Jg���-y�l��5��_���UxU��9M<�	�f��c�4���I�V�!V����`��"�B>ka�-������%LȬ�h�S`b51ӥ�y�7;�FZ\�
�#.�S��Q2�� Y�k�>���@�E�����__���}.���Z��{+�:��
!W���͙�(�r�Z�0�^J�����/\[P��h�lR?M�
ZB䑬9��8Y�ۚ��w}��E>�3����x�8�81��wQnn�i䷱u�����z޵�3�Bp�Z\��e�RP�0�tw���8�y�t���K����7 G����x����)�p��B�q� g�;������������Rg��7�w*�]��!���?��E	_��t���j|R���	��q^�6o��SΘm�5��r�(<M`�o�s�r�!�9&6��N����+�{Ƃ��K��N��Y��5�CfL��Θ�G������b��&��]������qO6��GƧ����e���U�ϕX\��>R���p�NW$M��T������>���ړ��L��@؅�d$���Δ�Ҥ:W\Y�4��m�v�|`�[�l�is��)��*�^�����+x���%<%g��{����D	v����Y��5!���Vk|>��c�?�q�J�I�q쩕�㶉%���������^�*a5h֨}u��)k�yc����0kv������ <�$-8�~��پ�9ލ@or�8�fCH*�l�]������`���1+L�xk��M��u�o����.����?���8��w��m��*.�k��	��[*�*R�������v���bv�Lm\�v�	��熥����wϖ�ֽ�gZ-�M&x��*�̹�9m�e�.Q��$��l4�Up<v�f�4ġ�"_F���-�)v֑2�C���/,��0�������zRy�ɩh�6'\5�U�V����IV��!��@�����l����Y$+��`�ݪ���{�(M��Ϙw�wk��ri
��~��K�����\���T�����v�cf����e`��D�\�5�I��z�������8�{�co,E]�<��o����S�X��]_%�_���$����D��f���̂�L�` ��?��з�����S\�d��n���ߛ� Y����*6h@/�{m�-!J��~�
5l����g�m��ւ�c�7��[|&���ה�isC^I���f���}�#�hHVr�1w��zgf�(Y����5uUf����K���q�K����u7n"�V��}y�y�}!�'��������4��p-wخq7ܬ�S��&އ]�UP�~
I���x�jC3�z'��y"9&�Lb��e�V]�]�

���$(l]Pm�ē*t����sw�ur���(+W���M��*|.KMQL�@H�ztw7R��j���mӹ��Uƹ+�K�|t
@��t ;��,'� �n��2ŬKZ�kL�=��th�L��\嶕tt������%[�������VnR,�'�q�)�̟���u(���b�/�����sr�U_K�(��~3*1�z�v��l��c�s����o�|6)�~a<�Z�F¤������0����Q��3����鷙ߪ�1�(���A~��B>�"�~2�[.onU���;~\ƭ���u�Ga��l)d8��ψ�I�Pۖt���\�3;����r���vb8m�7*����Bzi�>�4�Ĺ	�65����hZ�AZ�ڑ�#����ר��n�KJQ���/ú�1O�'F���!������ �781,��.y���F��:S�"(����8>�����''��-��3��Jv"	�k�ר�֗6�.Y�7�>/E�N�Cg�&��9)M�h����L��[e5���q����?�F! �<�g��c⡸c;>Nd|�:R��x��"�+Y
�	kƬ!�����k��n�޵����-�?�;�@�ԭ��k3�x�ѻ>��u����b"Ԩ?��q�3H:rݷ�upq��È�����x���u�`{��`���q�:���he��+�Ն�,u��c5�,��US*�Ō�=�r�0��L���љ�N�֮��/�o�"����� ^f�]�q�-f�tl���5�� CM��M�NET�Q��T|#c���@FN�|4�O7��QDDDp��gL���=��gޛ�I�ȵ"7a������%aI��2��O6���gغ����a;�U�9���Q̏If̋��|���n#�}�Fϰ�%W]��m,U\���׿�������mV@O[��é���g�����D��D�wEBӿ�/�`��A�G������K8PgS�(�}��)��..�Ws�^������[��s*��q.[�����	����ݮ�b�cB��Ҋ	�>6����]ە$���N�[�Ǽqm4�#0�S��Y�ed�44�rhY���*�"2;���	�Ф������Cea�}�aRO��a�0�F��:X?�s��R�?i^�9�����@
,{$�z������S��rDiހ(�D���50w����N%�hE2@g��2Эwa�!�n�wΟ/	eu�ܹ��_��O�+�cBvU���/��1ש�_�;�� ��<d���/����g�V���Xr���&���У�������M	�6D���.��ll0��C{�?竭b҅���G��-7:�4�?u����S�ɷ����HQ� ʄx�|Z&u$EY�TN}ϰ�CRB��]̬�ٵ|�&lw�vK�S�6�k�zʁ�r��1vG��eҘ!T��ӑ�ɞ3����Q=��!B�nZ��vZ~bL�ro�q�v]]]$����3���M^%��{X��v�������)���k���}/��z�G�Z�4fu�p���72�]��/ ��'�Xu#3�P�)/q7�6�"k*E5��/p���Gb���9�y'~IE}���:X���ڨ����;��X�W��f�p�ՙ{~rZIӷU�j��)�J51�;mo\o��R2�Y�{�xR�V�����d�YWiQ��vZ���F�]頃�UB)��ue�m���!ϚC!X9Z��3c�y�?;�r��;4���o�gN��ܔ2�T��?63���-uBu�����*��mG�����r���
��e6��)ϑٴ����ǂ�F����|���]8��%`K�%��ђ[�O�V���^'���8���w �J��Ȧ��3*��@�S������RD���� �˒6+u�����T@�%2�YC4\M��񢢖IJ��C��\��e5a��,q��]�{f������&=�����*\�/�1y������Nx�sVjZ�:2a"����A��ba���|����� � ��UQYp����r�������S���[�.2b1��;e�M��{q��z=ߟ�a�l��*��^^���׶Kx9Ԉ���W����$�������������KҶ���M+�����.��p:�&\o��e�?�����|1�?���A�|��(�ZP[��P#hځ�c_���ٌ���ռ��a+���ֲ�?��!<ɋU����D����Ђ��p˛����kt�a�ㆵʤ��R�,��H�	��Z��8����g)�)���JOx�P���n1��ف&�$)Vof6��+�A܎�?��|�P�2���ԋ+�n�Kˊ�^��/�_�j�}�S!'P!�Xϟp)�tw�Q��Cx�S�d�j$��i���㝺�h��N��� �Y������ۏ�m,�a.=��N<�XЌ0�54�}����{�L6�І�Q�^_M�\Z׿$|��;}��N�0C��,^͋�k�C zgW���5�)�j���fl-$Z3y�(tFT��k���!�h�2&{�9-2�����1'C�CE��u�|��gE��x2	"�J)���u��Ξ��;C�Y��{'|l={�,�������%7�Q�c#˽F�9cw���kɅR��/��!Rsoǹ�/�&ٳ��!\��X�#��f,z�s���/�Y���6�5u/:�[4�,�����E��-�.��d��e�J[�ߓ��܂^b��O������:y:���O�OgU�#���f���4��"�݂�|�|�7Vi���w.`6!߫�rl�m��賬�{�bI��"sB�y�hȆ$�?�����"(�޼TBA]`�X��/���,b�	=�:iq5���c��hږ I���y^� ��)�}�^���?���L^��zv0�z�DN�<{9vv��Y���u�aP�ƀ���tdѝ�1��ތ5�(\��?�h�C3g�sM�$��C?a���
��|��hG����{߿
���������w�w�fo7�<�U��d=~�r�V6�i�� �V�c�j�^#�#�C�
�ʑeJ2�r&����n���1�'`��z,]��A�a���5ݜs^U-|_�G��b�p��y)��l�4�&�B2�iQ����9}!pS���O��=�Q���Xn�D��,��o�z�[�]TRs>����z��/U�����+ދ�>�������ן�8�ޙIƸPK,�3P�#�1�m�i��=?�H���"�lXC�O��R�x��8�����v�_���<���:<I-��2J��^e�(�O:a��;$8�:�p�:h�+��<o�C:f�,���:W��;a�t]I#���A��{C�/��й\mnY"��0w[: ?�s}�9�,����.J/	����%����ӵ0\��WN״��ǿ�^q�6;D��Y���/�9����>q�R�����y�UJl9[���R�B�L��X�~%o�Pgi�t���;{Є	�O%nud�ʲdn��6iC'�c/��n��g�&^}_������8�/&���(X�����2�H�Ȼ\�O)����y�1y�|���C"��eq�L�5S�������.�����?yx�Qq���h��d�Ui6p]N�mQd��o_1z����+�vYJ�0�u�[�i����6<)���G�2v���� ��`2O�ڃ���bÎW� �F�y��&�t��DP��c��Q~2�rDkb�͞^gy�Г4Ѝ�*���'�[�"�����G�����@=���܌��D��6uT�����z�v��W�>��_�$���IY�_�~�P���>`�u�p\����&�v����%ܶÇw .�|̃9�~�cBw��U6|�,�a��ئXWx�f���(��>݄�gOl�c�wO����ݮ�&QaEY�l�!��k��?[u+O�A����Vv���%C��Y���'���1AA���^$%{�W`���sR� 6���hpm���H�m:����j�-�j��?���dz�;�#��|�j��ZAp�!�FB���z��3�
�
ae��fUb�z9�b������S�cd!ۛ`���<�v��=��g�#�.�n�f[�OΙ7u�G�f�.��#x��=��������&�*�+ⴠa�opa�,Kp�E��m��ߴr<��8r r�SY�\��tn�����7��v�@���~�_�4�����֊<���3̒��WPN��'1c4
1��TҎP�Vf�]��o�'-;�gw�p�с��|��_�nY�}0~hRme����ѴHڢ�4� �ǭ0~{H��/�|1a�X/��(��T�I�s � �
1?�k=04i@����]~ƚ�n�,y۾/t�V�f6�.<��_a������-�z2��5���SI�Zx�z���L%�0Zx��%��F<���;��9���� ĩq��J=P:K�$�|V�b��z�6v}%�ni���X '�~Bp�.��'{��e.ᡝ��{|���e��e)3�x��SY����HWb�u^*��|mJ/��ǣ빅�53T��cc"�Y�RQ�!�0��t�!�-��<b�"�]0��_.�9��^�֯'��$c�^�u$��)l?�IN�5�?��.M�S-��ȣ7��Y�H(��9�01���M��:	�c�����%��Ҙ�h������a=� �[��߽l}%f�(kF�q��P�hq��f{. �M��d��"|- �/�k���-Ccq����(h���W�A����`(Pvu-B�a�k�Hxۻx 	_��+<2B��ٿХ���"G,������>��n�k�ׄ�*�ί�0���U�0�dwz�BH�?�-j#��rr���/�C���}�&{�㵡c;hB�	��tȣ���0a���\f�L�܎�Ƈf�A:�=;=3�������>�4�9�.fgl"�f�x��賛o�ۙ�F�~��-J��F�>�6	���T�����B�4n<$�_=+YF��\GxN�L����pUPЁ����p�����>~�8|�j�,L���~�^aS4YƆ�����'�֡�Dg��3�WHX�^����Y3�[n��1�"n#+�Z��׎��H�(��d�dYfb��2	��&��u���Ls�i��1)Vzd�2�s��d��/�>͸ل���r�0��z�������������F�9�5P�~ʟ%&��{р�{�Ӣ�˥}��~�4�u�8tI�U$����~�m+�-�� òh�/�<.1)���JT���L�P��|gRAv����m���"�m:x.l�B$b4:��t��x^�K�	q��]>�Z颎�/w�g����̩U)���Ƨ#�U�17R��Loj��/mz��YG�������\/�N.����ӻ۝����K������zOd������￉�%�M}�Q�p�O/�k�����A��u�6o�g����~T�a�N�VI�b��"�Od;�Ϯ� �w�A�G��d�����/��ߠ�F2IA{��V�2�n���jtzU�{8*�2������iK�%J}���{2�{g�#�@u܋�/�'���)s���d-����.����V�д�����ZM�9!<:P��t�>=�w'����A��P�� �D����R���d�k�
��31�ܸ7�"c�/�G��TbĬ*m^�R�}y^��LL��f�'K�И�94�P��"�\��j�O�_�>��a��tbJƄ� ��Ij7�t��@�ko;�pZ٢�6�*56$�����*�U5�|�O�o���5��m\���<��s�5��n�?2�Ni����EG��h}�|�����3�)A�/Q���Ң>���6 �l�tx�1$�}������c��IsL&H�A�"Hj��5�7&��o7J;.��;q���M�2ǧ��{�USB��'�O�)� �L�Љs�ۓ7�I�����d=�.�d�����5�c����ِc��c�7�8�Kē8�\}�����s�ګdA5`���8�c?���>�cxJ�s�6��e"�_�$��ޕ����Q�Z
8u��Z�'-��J�#z{%S*�0����M���ӕ�/�6�4wuf�툦s@)I��/�{�	�)�z2�S�j�^��d��\~��A: ��$ʺ��׹��tX���l ~�]��\�}F� �ǚt��6�;�V�xED��8%��g(�Y�Puul�S�������&8�ݜm�2�0�N�vm"�V,���r�L��u��]�Ѿ�&�\�ox�O���Vj_�|k����$	'E[�$���@<�E� ��8���H6ϕBl==���O ���I+[�LAG���s�=��;��R�	p�f\���_�k4a����bu����M��6}~M<Zo��T *L����ex���gT|<+&�v���-��(��0n���$����W��"%�'1~I��bB�ܑ��/Jb�N/h�ܭ��˿�uzˊ�uS�!0qh�i&f�"N��=��5H��K��6a��B��=����u�I�͐!��X8N�p�ȳy���!ȋ�Ȅ �
)44�&?�c���z����+�7��.�y�c�x�� ��j�����H���5vu�t��0\��\�5�_p�,4U�l�P��t
���(Y�1��{��C�S�Ab�G��5{���͑�1�r���$�'Lں$�b��s�v�a���H{y��/7R3�k���ٸ���>R,a�M�8#un�D�Ӳ)ta�-, 9�:0�����U\ܧ�:��C%���M?�$M\?i����u�˛�{wD܇-���C����giX������v�Mޑ�GC�����2%�W��m�G��XnaGiޚI&�b��2^vE&�P�r�dn�A��":�u�gJ�f���q	���q��.~��fQ���ĲTZ�r��e.Ј�LB�e��Tv�C���7��ں0���|=��s���.�.$E��T��z��vӕ~�����q�=��A��v1E��[�g��\�&�̐6	F�_���Y�Bs4{/"|�x+5��R��*�!B�4�Q��l1aP�s�>@<�����^S�gS˔�TH�cD,�'�ٙ��^��ۿ�r/;�?v%	�a��Ļ��t_�z�^�E�%����+��\��'�
1�JN�R�����Ј���o���yqWG�&� �ԥL��)7[�g���P9�k���'�ع]��6R��H؀:\VD��s�` �[D+�+ށxc_:.^�jAPƅ��$��*h܁,{� Us�W�u�-�V�~�!q����G�N��{�9	h���u�ϕW*��YHrH�m�PU�I2�}���^6��m�9��T/!����o��=�0���bb7C�����j�� u��lO�3\!��M� O3uu\g����d _��O�P
��40���&���9B�P ��w����㦃���R�|{�^Ts�qb�CF�B%z�_h��1R6�O������OH��3g���1]WPx�n�JLsH����Bs��[��/~��X ]�L��<� �0^��vk����[�3��(���R��E��}^VCYi����c����N��I�(���`߬'eX�FB������m�sm��*��ݟ+�Cʃ��uSG����S��q���_�L{�����ڸ�["�ڤg�=½=��~�Ed���J�/i�ArT�_�Z34Dθ��:e��8w,ͬj�AN��p�_.�Q�㊾6q�,s9����}�>�
KOW��v C��*Ѫ�Z1"p�KK����Xz|v�����A(qݒ���T����o" ,����r�;���$$R�T��4� o��IxD�u�2�Um��ԗX+���������fP(S�)�e=�:�P�sqK��K��vO\*���#�k>�(�X X�h�?=|��O���\<��ת8����М��.�D��fV=CS����e[��e�ӡ�	���j���b��y��[�MD2V�^�����yS��-�R�V�oS�jD$���R������q�s��	�ԉ���:0.��b�\�OK�9�Z��ؖ��'�F�R���N4}�RtS�d�.tiGS����~��v�Jf��=s;��!Y/o[�����=�l���n�C7�W#V���U��Rn�l�W�+e���(1���2�ٕw9��"���V�V%1��!ʯԚ�k�A:�%j�g��J3w�@����a�5��ް1�2/�1���g�ʹ�.�KLKl�drKg1�`詸TL�D5�M��᫺��&D�&�m�g���뜀(���L�4QJ:;!���|�F��6k�d���IF閂H �'R�p��;�#ƪD�����6#7Z67��l68�y�\��F��Y[�~W��l�)<�V�9c��3}IL�w��R��� b^"pfs���Ȳ(�j~7��XѠ7OkRydP��F-����g��Z�	��<�K+_��s��av��3'6��X-���c&�ٺ�o����ς���������'��y�\�@h5��Gp.>����lO-W諴~	A.TMWπ9M��Q�yU
�%������N�+S�g�	��$s=FH@~���(+P5���8��|U���?�_*�0n�����8$�����-@��$��@S�����}�e��ˠD;ٴ턄-{�����1��M��GtK �U��%����h�
I�M�u�\d'���3Z*`C�܁T�j�%�&��܇��Yf���;�9.$oE����gR<-�}���b���W �c*(�rE�zH�r7�팍�"y�`��,���%/���I��:zv���r���?$2�6c���h�w��=
���~|'�'P�9<��]�.�O�}7�|}����̄�v"���Y�LO�J��i�����b��lL��۰�NH/�MH�GW�>�{#�G�| �;V��.��BqA��Ͳ.\��B�%9�����*f4�8�8�!3�V���p�ӧ��HHrkI�2������҂�NCۛ_w��xW6�$�3$v�ǩ��֤�bq�%!1ŽWw���Sc��� ��n�G�#veDl�縋��P��2�/ӝ*���EQ���TH *Q���C��
�XL���@QI35)�q��,���,v���C�:����Ͽ��܃��`����8p�+�tsm�f��b֦j�D�&lS��'K��MU�ޅ�rUWk�5m&��4��-9즾�oι�H�Lzh߮�E���K���CPVu�z�JG��F4�a����,q�����'�צX=�d�?�OvCY������8ֳ�6��e�~�n��A�����M���>��v���啊��SHy�Z�̈���C��!�g�KT�<%����(��I1Զ�o����˸!�4D�f�):0�(�b�*��W(C��9��f[5��J1�p�Q��Ыk���JZ��]�g2ޚF=�<���ް��4���Eڈ��'��7{��w�D�O~���x�M[��0�囩`�>�+��"�c>W�2�v�c�k��3�J��Y�� D���Q��  �ާĦ}��\��m6�`Ӽ�V^� �1�D�g�ȳȦ��+<x�(���N���W�gKR,0�d�멏���r�mP����q��.C�z�hX{3Q!R�Ik�-�<��`��Ξ�>W��5ڤ�:��˥+��U:���pħGj&;$�#^���I��^+Nr'�����Bu������o"X[x�h�iu�8̒b�eBu.�^I�k���?[h����J0�o:��h�:D;@�S �k�9�Ci5U^�D�ӻ����R�qɆ����ܽ7��\[��a��E�^<�Rj�.�u7pٌYV���mL?�z���aw�{J%Y��_��;?f�����@˧�+���uF1O����|�g!:-X���2ESr~a����.s1Ze�k�ͬuC�^�&l���+�^���Z�X]�<���D`�X^��ћbw��{�$s��9 M�xAD��~��(���)�QJ����o�
�Ǹ0����>d�E�W8�7M��#��2idq18�)�k��(��x������V: �0 4tC\�
e9R'�{I2X��"��𑠗.���"
1�a%���Lt�/P8���p�w��@N���n(ԍ��5�ڞ0�z���3	�$D�����4���Q��҃��o���w3kC�Ó����6S����jJF/�A�ɞF��=\K�Gn�G�"%�W^Gb���]<�W ���lP��F�zs��bi��e8V~��Jt��y(����p��l�t��+���Ѷ�_�k�IS&O�� �uȦ�I{��2�Nj��LS��+���W�q�\G�J��I��99�6�{�C79��&|����������/Q�9ċԂ�!Z)m�/K�xe�8Q�%��%ҺĹ�!Wx�ʴ�
8��J�=���%���h(K(��2,J�Z������\K��4���_},u/VV��!	�G�ͬ�����8] ��f�e(��P76d�Z' R[PҪ�D�X�J'�KA�\w*���+�\�@�l�\�SϻZ�/�8b;���Y���?�����,��(�R*K�6\�79�m�Glv$i!�����5�bȿ�(��GKD�{�UQ>�1Gl����<�z�"k'����i����p%NP���j���dL�RG���[�(�oXֳ�����`�6�>��V�l*m����D��J7��2�ye
X6:L	��J;=-�b��E�'����}�t�/M F����2��z�8'�Y1w5+�\����F�|G�N�"ҩB��f*�o ��P?�/�,;y@����Vڡx�V�.�]�ZY�G���^�#P�F�pL�$oI�;Mq� eɚ>6�s�跞���B?D����@\	����P��V�Bօ;&
��8|�T�?.r��o�j�m���4N�&��R��νHO� �
7��*X�lN=�
<���'�z�
�^��$w��Sˋ��D]ڼ��P��?�,Gm�;�0��-� ;��(<Ѩ�aL�J[���^��᫳*"z'�9am�.<i��l�o&x�;s@��{X-�6G,h�}w���d���Y�O�(D��fd��v-��1����!'}�P�ۂ�2W���s4�C+"PB��Y_�`i_"}Tv5I�@<���=J%��b^F`�R��dQr�Ĭ�U��^�5�r��]IW�S���v�I��{�� &��8����v�*cD��00� T(��X>@a3�v4#���KU�<��/u�����i4��"�3&��Dm���[i�g�ތ��G��3��i0
��7L�)�М���y�!��\��Z]i��b�����v׎��ܶ���C}X�:�^N�&3�@��uawyƅ�M�*��(w�]2��YTP$+��cΖ������\������]���	V@9t���eĿ���I%�RD!���>҃����?���V��>T���vT�R����0t���#��aj��X-b��8C��X�<W�}�n� A>+�Ysj��m�Uz��$ҡa�a����l��vh`з�����X�K���u�W6
&���y���M1x�.
�� (iQh8����D%i�lxi�L�n��6qy�n��^o�<�a�qA%	�
`�e~�����:�BN�K�NP4�����^�>�EӾR�ajL�s�����S4q�Bs�&�~�g��^�<�K�T���s�/�r�����aQ��0��3M�Y�^�e;��F��v[�^���Ox���q�s�l�}�4W�/�>0�p�d����2�@r���vO(4�
�|%�mdm\�;���Ck&�z��K�55�w��]�5�AP��`���7 ަ��E.�)y%Z����Q�Ʉ]oH�h%�D<3ŉU3��<O:��C�h���3�.aJw��z�s�����<٣DpLQ}���B�k٨���+W��������y�.� �q���<)�a+�y�dC�S#V�l8� �i��To9:N	l_���_�����4S� Q������1f��ex��%ۭ	��{�IXN/��1�q�"U�E�e��˚yc"�uZJ9'h��a���x3��۔�aG�L� ��ױբ�1�[Է;D���;*C��2�WUk-fM�#U��'��:H��w:�5��29���z�%�(����dSݦ��%�%z��n��� ���6�n�dufL�	�X�?gl�O��V3E?[������4/3��:<0,�l�ʞ�/�@�NP�I�-ul�L^��=dS�Z1�to"/��)����:G1��	&Yd?��bGA����8!z)
�Ue�8�%�9#��^��Qu���Q)����/~��	A!�DN�W�bk-.�[ΑX���j�&���h�E*Ќ�W��ѦG�ĵd�	���%B�D(�O�����r\�����I��%�K�RF�*�m��b��.,h�i��MJD
4�䎴V'�mp�=<b��wP�Jw����?�l1�ķ����3�?d�9kaT
	յ~P W�ɶ�ȓ d�� It������.I��3y&2"�v2�]g������M9�L��q�!=P��8bK��O.�����d�C^�o�60� ']�P��W�WI3ީҐ�mg ^��J��[�r�3ڽ��kd(��o|�$��}%F[�1��:'��^�$S:���}��@�^Y���������&�x桅��r�T��	mDI�J������nhiw��	���9ίJe�x��ퟺ��p^F6l�b��beS '�щ������?Y,�M�4���j��
00�v5�p1�����R�։�������ҥ���@�s�Tzi6�g��b��+���ήf��;��$-,�c*�޻,�]��v��%����B�h;�c��lp��ݗ t�z�R��k����Ab4Y��I	d_��^ﰱ���F�
�n���	�8������.!��g_I��\�Z���2� ���)Cwō�*\G�.)�ֻ��k���o�GF�D:Y��ը���Ȩ�BNm��Qye���)ۯ��U�P�%қ���u���-a�,�2J.�1�:��p�m�K萲�x��F\?|��L���j"����"��6Ľ7���皎��_��}[��t��M<ν$u�����ZnrHY�/=F�k"b{%QF�&\�y���Ɉt���+�a�^���"�@���כ���vX<�����<�����K;d�@�oY��<i�W((!��$���6��I"l�b�?��g��j1��\F�"��$~�#���O=K�5�ѽ%kV�iޟ��Y����z�ϫBE�jO|��$���X�S\OM6�^�Ĺ���?����r��4��_���RK�� OO3PB�d� �|m��~��#��#(IP���ܯq�FfB��'�l�cAf��)�_�9�2�Пi���6��YZ�@�g�������+�ӕwj�'�h�7\��;�3��Cv�+)f)��TBP	R���$ϭ2�t�MUV`�#�+	��)�T���/�ȹt.?,h�L�p�Z�A�L�'Dǝ�}c���+��j�*�w�DH�Z{R3�_�Tl��o���ʡ]Y_,�5E�~E,3�2���������n7W�Dw�/�0謾��"t,8B�S;��m�z�ys�M^)�5�E��M�4�/S��^<8a���pE�Z�֭.%�ac�;:�U�
���C�ZYH��Q�Rp�i^��H�1Z����֖.u���C�ˮ_Y�ב��f�+m<[���Ԇ��lk��u��K�$(��Ї�M�		�����Z��d�@2��W�TYt�W
FhxΘ�8�Ui��#����؎շZ���i�-�1D����sZ1ąm&46�g(�WkiWU��hA�N�}��x}��@���cD�����j~�].��vzL�5y�礪 ��Ǘ��H[ۀ�o�pFYG˶ėrn:^�lY&���Oj��?��!N�t�[��N����p��w�������K��]��D>�!��#jX�&���V!w�����\$�Tm���B�U�G��D�|q�k�C�j-J�%-m�W�#�k��~���H�_Q19�-�%Z9.0~�G�YQ��*8ME\��"����Q��b�C�I�q���+�Ͷkt:�ǿ���c	S��� �_���#�'�Y�B���Q<_�.IihƼZ:�i4O�E�-�-�okp��[A�/a���)~X���z�7����^�^{?����V`E2-�ۣ	�C�����,���ղв�#���+��� ����Mf�\��a�o�{�F9[Uir�4�Md�����A��*���\ӱ'FB�2�_�S�z��PF�&�O�������g8�L&��"T<���Ys��9�P$D���ANf���bk�Y��6�l�e�;�Qz+�Q;�4���@��0y��G�\V۠�JK����݉ɻ���Բr�&L{/R}K��b����T�ԕ��"�l���?2�N�>�(�������|�汉M0�D�\<���HF����*������C��'�y?�3�ѴQ�ho�㵁�n"J� ���W�����T��=�꙼��a�}�s��ى�e6���ӕ�$l����Nh&وF�fz����L%&k��6?�sgHg�	9˴��WE0�l����t��/=��A��i��n��y�dB��1i�(�9�����Fq�Z����zӾ���!W���w݆D�3nA�,�
�R�n��^��\k��t�1n2(�r-�����Roqy�R�gO�mk�!�N�Qn��n�ٳe�_�<�
5�T�������=P�'^��(k_�m�l�ƐU�� �
S��i\Yt���K�&�L�:v�/�B�4k��}��a������L��B�R׺�q�B���n�J��џrŠj]ؒ�k�g�r����*��ﶡڶ1��+\�@�����*�V��.A��f(E����f�BB�DA�{i	��f(	�zh�A�繾���̟9��^{����O��wt��И*�wT~���?%)ģ�<��m����o�&s�_p�:w��"���)����Uq�|��'�;����Lm;�ģg}��g�t������(��3�+�P̞����9IX�8���t�![��r���/BK���U̥B�0�!�����/�_�k���l�zVZ����=�Ŗ�NV�I퍊\Nò���H�,�;>{�(�������\�����˜S�?|9���ч���lR��lz|��TWd�'���SF��E��$�N�`��w�X�ٲ��h�ڼ������[G�o�U-���	���p����b&��	��������է��X���@YC86��o9�=rټV{�'%�Е���Gw��'V-ƃO%wU�z�c$�~��?Ir�4��>����<��&�:T� n��&�Y��~h�'m�ѡ�_����8n*7����B�ê����2w�E�J�3?���e6m��Ӈ��f�N�X��ֹ��~�a�p�:��%�<�%]�D2��gb�2���I�(�[�O�o-A�m���=������ܻ�2�2���UR��?��{�I�<b]f�43+|��2�@h	�q˽��uV�!k����2���G�+N�{i�I��s�w8	:T�Z�#���r@q4y�u+���Ƅߵ>�SWu��䌜�n����t�I�;�vX�U+�ǂv�q-�agQ�L9|O�c���_ͱ�t��Q��)����F�-1��U�ڴ<�s�$T^SO1�K���&Fu��&��6��|W�}�P2�D9{V��,�f���߇w�2�2�C*�p׳^w%���,���P sUw�.);���)j�4~�t��T@Xk���Fm��0�b�����S��q�3.�ذ�M䧅�%1���"���eݾ
�T�籇���n��_��ȚR!$h��xD�lZX�	t��7L�oӬ�:�>����U��������@�՚�x�=o����ۀA�f�ӌ��C,FZ�Le��?��["\V'��	��uS�3ȔI�RS����I�ՑO	}����ɑ���³�0����C�r�%C�Ig�-[p�˵��O��)�_����U�uݪ%��
��HT�Y96|g���Ǖl�����XR%���QhA�gL�T�$D�@T�MۍȊ���=DM6�~2���/�X�Y`ʊ��	��!w)΢�[1�u��NU��I/6_�қITY׈�8��ÚT��N�ea�u�ę/�����̀��$�sF���5�)���T6���w���#������z�z<R��#�*J��靸�ǜ�����|;�6��L�_Z�YL��@26̔կw��������S{(s�žT]��{���>�j���d��D�������/�u���p{+�)��w��jn���P�^���V�������<�M����
� ���]bskQ�4Ro����u��Y��A�aj���л�5�]∇�{�FB�+1_��pp�c�c'/,�+�o	&u��^���Yʻ@=��F0<Et��J��YYI��|c��S]K3o�:��	|��֎
���ur��X�9�D0�ԃ�K���-�/q���,-�A�z�6HA
�I ����$8K�� n�n�rleI��}��_,k��U��J"�6�х>��S�a��?�)��B=�J�zVNY��cf��5��v��3�b?��Cc#ļ0HqI��L�Y�vE�N����3���ݗR��uɁ�?j&��Q]T��,^�r���v|%�\�>�о�!z���7�*�%n�gn��|�'�J(�ɛ#2���#k�{i��$p�\�ȅ���X�@�T'����l��O霈��YڰJ)��H�bOBU|��^���d�<S�vZ�K �m�q�A��u�`����C{�s^��H���N".o���b�	���+y>2o!�٦��~C���Hl��K��:;�LU�Y�[��yg�귎�;DsPM�n��D���#/��/��ۍ��=.�����?�)3S�7�3I�����k�j�xP��W�}��i�;�#��{�]�D���+�Y$���6�GWa�z���
+�����z�Ё��߹ߊ�X���_�ˌ�����f��UT҉5;T��f?RmJi�kx��/@d�r��Z�"r�z�)�U�Q�o���M_O�޲�Gk��8�^���q�C��.`oeŗ	�R3A�%'̫��d�IU�����[���ɚ���S�A�9l1*÷�Ҋ8ف�{tf���*���n���q~�:k���

H���4�&i�4�׭�~�5��-�z���.���60�'������w�45B�
�n��C{	 ���������So8��n���e9��������O�5և�ǣ3ر��7�����[��	��K���;�*�q5	�\z�j
�3��R�8��Wh]DzM�����"���8Lc�����@U����^,C:,8���$��N��*)G�j�.�4|v� �N-?�r��5r��l���[M@�E�'{[��ɾ�U�@�G��8����E���G��8���G��YQQ�� ܛB
M�/�d��V
���=d�%?
jYw|AQ�->�R��ƏU����^�Y��g|��Σx܌Zޭ�и�؟+�t@�K������m�Z|�]�
��H)����:�\�B��������v�]\k�����iʆ���-�:.kT��YX�m��*��0g���$M����2�T+��S^�&���w@��L���K9��bV��w_�j�AthH��
��uȨ/?S�S�������Ϭo�ǃsk��(�1�-�X�:�p�4/��9�<?�R�j�AD����`yS,˘}���8:����%��>���(�#�fV��).�������nN�8-D�$܏O��H����+���E4��>"�5���0V�|�r����/ٲֹ��+���a�IE98#Ut]�f�2ܣ,�ʻ��ړ)����5����0�����`*2_�`7C�]m<e���F�µ��}�p� T�y�O�1U��:ݑp?�[�_e���{�շ��M�}m<"�NG�>��I��6\�c��� �
�]r� ��e�����iE�Ʀ�gJUiEnj��R��0?��  ��ef������jK���I��#$������p� ;��X~&@8˜�1#J�fMÀȱ�V�t��	��(g�XY#����7�g�E�9ծֲ�Ψ&�����=�u̲��SNK��Y��Eɸ���R���+��M�c�z�,}�zY�W�Cy->�l�Ya��AK��"O�̦8U���X�>�Qm�%�m�<� �x�?H�]f�3O ��d��hr� Ex�]��*��Ƃr�Q�۹+ �K1�'��&=K&6���l�O!����������]��]��s't�<\�5���q�^EXҖ�)���<⧼ �	T���~��.: �q�I����S�C�ڊ�_Ǽ��ʆ�ѓ7�ZsT�'�.�3	��	�&E�rE�o�nfPl��5�c��uVz��(kR�W�t��ɡm�qIx|�q	�������=x����5D�~ sAiU��b����Q��JC��J�[f�ZAx���|�	�+$l�dW�/f�����!.��5��ˎ�~�W�0����6[/>�]�{d�7]Q}l�ܺ�1����{��Զ�Z�ﭻZ9�yAݾ�F-0������!���:����t�oZ8����������Fi4L��~��:a���Jv/�Ip��UEҌ��;�7kگ�B��m�=mV����Z����k36��W�	oXg��i��?��%�b�
�i�bf�t�1h�C����ަ�uܳ�������ț� ?ǲzV�o\eǩ���ٛ䀠��:~~�����k�&=8B���E�ԩ�=K�SwUJ{��7
=:�������5M���I˛ym~�w���f
;̬W�l��}8$-Z����N=����?秘�Y����V���_'j��C��8����ZM5���#}��z��oa�r�W<�r3<<�����eHxp�8�>:�o����z�^F�7��E��}�2bbb[����V�����m��~��G�}�":�^��թ�杪��"HZ�4V�4��'>����n;L����:����!55�]�M����:eK�szr��;��B��a�a�m�O�@HC�]��0��b�����O��4��L�)I�[k�;����qDh��pD�Tk�_�ߴ�J�,ڊ%������rd�{��pf���z�
"��5�&o �AS�/bߘ=㖙b~���bs�`�6w�i;fi����(���߽u0+xC��
}��Q�a�R�J84+��A��.<���z1��c�ώ�>��Q�x�<|�a^#�h��6�w,���y��@#��yF,~�<�QʿL]�?a��c�;и71���"�20Z�K ł/�q��,}�W���Xh�{��?	�*(X�Zp��so��#wN���ޤk�)\�!$inl|ӝ�o�����`�ֳ@/��y�>�q�'�������݈�O|���	�4�<�X�A�u	p�"���O�x���k��1 �)#0�{��a$�z���e�U���D�,)ÿ�2z������)Q���7�"�?����f��\���>�ٞ�^�sQY�>���ӕk�]���R[M�a��WNT1��$0�U/qF��8ٰ�.��b�HA�A��_�jVv���<n,czP/µ�����(K�s�/�����V'�P�nڋ|��}<F֞�ڵ���og�P޶K�g$Yo����6,.U�w����	h�pcf�ψ��,���I�b�_�>m����ʻg�PC3O����7�{,c'c/�MbSa���ċ6��{c���Ɔ�Y+%�"�i}iR�X�z[yŻƟ���a>��)�iD���9�^w�[�8QIg�ŧ'F��Ws��Y��],�bB�cHF��b��/���|M��g�S�Svs��M:n&* �7��t˱��fS|���~LQtho�Y`Q$!����a�2YN��'�(v/"]-��]�0nW���_��b�@ب�����*��"�zNuU�մ�g`��:6�7���'U%����م~�zP�[voG�x�l�_�U��R3=��� '�ki�1%�Y����:rꋾ'��}8�	ˊ;��шE���Pس?���7��3x���I���>���y���tQ��"��K� ~�.1��4���5J���?��³����J�`$lvil���"B�ǳ�Om�-b��ʁ�ZIY���y���Vn�����i��;o;��=�z�t��u�d;6�I�-zj����M�݁�@�7�<A�^����o�E�U��baY���#_Bmj}S�R���u��Z6����7NW���z���b2k��B^M�����_�k�PP�A�Db|�19�A\�E��J�n�Ix�W4�/>C~�-	9�_�Jɔ�X�B�MѸ�=+�����t�u�������z���4�-�{p�ML���G�,'Ye����[��K��|�$�={Z��%�ny��hY����R2?K\r@�7U�����E��ƐE���
�t|q�����p���O�*z���0��z�Tt���@X��%��'rߤ;��[��5�y���^���=������l3�W���5�̓_�8�w6��/C$�yE����;k,BX��e�|��0�X<�T|�>�?�	�x��I�Q%���7j8���|�m��K��5������c��WG;VY�AIͥ��j�Lש�q��,3iM�SA�a^#��R�UJ_�4Q���7��K�b\�Oc���>L�����g���'(�H5f���W�)d�߄�w�ȵ��7�Z��B������f��0��`4�ܕ������;�([U�=��<�1����l���3]���g{�5�F�i���oթ���g<N��X��P�%���.���A��b��hвq�,���?��Ԭw�j���n5�ԑ�+�\�>?����|�u�t�J����U��G}.�N� `yZ��O�Q��~S�}�g��dF��`�4�Eg��Z��Iډ,�,�U*� ͫ<5X�A4P��>|) �|���>/����R~d�eDC��@ͬ{(�
�>�ZT�.º֞��-.��ao�m@3�����0��X�@w�7Ҭ���`���5:�y�N^"f̼�V���Xȹ���p�[���x������΋-!#wa�e}���]�>�z�iÐ�N�n��1�t��"%��~��u�wb�̫���r��5�7�Z���Q(����%CCjum�����Z�h9	��AGR�Whp��u�2�8B|γb�o<���,��7y�0�� �a 4�d')�;�u�J�����r�[���8�v�Ƙ�l&���=L�R��!#Ѡ��O���Gm�ҺN�����%L��Z�RoYo��r�\����(U��kk���Q0��=4Vv��D�U��0/�!RN>3NJY�h�2-]���i�����W��0V�<�a����7j5��&"��R��j�)��s6��=��~{9����8R�A���e�ݘ��Le�N���0�C��&D4۟:���e�D�ay��Dk)(�X�gj*�Vz�ů�f�t(/~#8j��C�'�E	)��2�M+�ҭ��x��z������֣;�����*�H�V�J���4�~ 渘����w��9����R��h���Z�F��&,cdc;
��Pl��2��\H=�#��i�A�`~/ ��s�|����Se=w������v����[�J�.�č�}HI�tKj��Z����2I�p��ZvW�TN]�n�Ā����/�̛9m�؉D�XՔL9�<�o�0���:uN�}�U7�i���',Pl�_MM,SU��)Z����y@��\��/����"y�-���(���y�P�~́yu� �R<�ԀO@�u�a9沦#��Td>��{ݳST�8����>/�S/,�>ƫ�"���٘!�4��
��4���p��>En�bP�B,�у=��g|�*�9ۋ��&��/�B:����:m|�C2d���l��i9؍��	G���_�<���b��փ����1���i�P��%�ǥs��;�q�M��*�K�4�5�֒ͺZ�Cɻ�}�����Y=u��8{g4�)��~�e�mVf�g��Ҙ�Uf�(��}h�^R)�����M&G�$��m����=�ܨ�{��bT�O&�w���t�ޫ���!��÷3[�X9����E� 2��z4�s���.7��4?o��+o&�7*�8dF��+c?��I�}���A.u��p���������{�?8�È���疠?�7��f{<W���9�5��*b�i�WQ�������o�!K�V����`��
x����G0������vd���楶b"J��]���J26�A92½���C7����n6�d6Ms��)@ZK$C�ᕈ^��5�w"γi��ח�1x7_ '�ZOa�y�}+3�!���7v��r�	���=�$e���e}l=$�?�Y�����\�=��l���zf_��*b-�6�Q��q�Ѻ�n�9�2b���Lc����礓
W�F�c�$�9l�
u|�.��]R{��q|W"/)���}���.T	ٳ��#�T\��1x�4='��w�AG:{'RW-Z@�v +�j5����x���2��l��e��Y�; �bnrHu�Uv���i�
��<v;;;s���18�M2;�[�{|��2%/�U�C���-�
H��f�.�M�'.8WE�uQ7��o��2C9��gIm�~|kj�԰I�hg�75�Yyxŗ�c�*g�nw��}�9m���Y����83OXG��008� �푴A���~PY�C=�u�����_�#5�yp�}�I�� ��w ��O{�����r�_��!�hʯ�l�-����qoڪHp�"zt�̴�6Mr�e�D���2J�I�	�N����j?*���� (����a��?/�d�$�3g�02�Z��b��?��mJq�}����^����#��c2��P�h�u�qq����oE��a���W"j���ǑI��-U��K�[��O��	�ond�O�&29F	�w'ܴ
�%#�+�^���ӜIi��Ȟg�~�f	��M�T�~뗩��{ g�I>�@-�B�X�߀���o�ا�븿�n?�0L`����yϠ!���q�,P될q���3Q �����F�p߈қdK��.xNA���U�aY�Ӊ�7��w�䯫C�����i
��� u&!+�1�i�F��k�Mv �[�:�IbTT������$���ƧjV%����s��aJ��0ޢ��T��"�X�J����]�k���ˑ��b��+��=j-�,;m3���-#��[�*BS�4E�L��J�n=?��p�l�����o�����p�^d�j��
ӏ�b+kk>��'9�;�
8T	��~���2�-wT���46�p�y��4�ֆa�U�6>Rs� ��y�L���F�K��}TF�c��*��$4�_���s5m]���R��c
�>�E��: �J!�:���t�2���4�.�[��mlX�.�giߞ=-G1���6�-�U�Zco/K�+�o2H%2d���u���}����eӥ�i�%���e�H�U�<m�Ư��S��ъJ�f�ce^�?��8��t^��p��0���n$�}`ո�ʣ�T�5 Bd��:�ף���
�{7y�i'��@u��)��X�	�Z�u{�й���F�ۆ����ޡ�̿6�1X�k�KH�JH�N]�<VId~�
�
�2VϾ[�h�?��g򑼅�{yF�L��D�'d`iŀ[M�n&G�#k)�e�K������f�/��=�=�d���3��>�%X����
~f晋]�ӊҲGS����~A�H���<1�I� A����������BDB��k��%*���]Լ�[7�Q��X�i ��whi�g������g�0�C���"��]�f���2���*>ˇߌ�y��.I�T��f,�U����Oߎ�Z�W1�06�\n(e��셔R��du��1N�嶫���h���G}��X��w��q�����~�l��� {���l�5[��ہDv�Az�OnZ�f���;��W�
D���ׯ�"�2O��)~*��3�U@���|����KK��I��È��
lʫ� ��	�S��h�+�Q�X�h���$!A��&� 0��3��vY���=rN:����u+:*wY�����Q�~�I�KxE�EdݑN�ܯ���>!������#�+�q����&��oԹ�T/��1�w�����_�Ft�D^����2Y�����6�9j����%hRH	Rތh��A�/�`ۛ�ra��ZG�����=г��ExM<�y��=\����؇��%�$��w�N��d�u���ۄ{PN��b���+����Ne���
�x�{��r����}]���Ayd��?�sh�������L�\1�yL��[Sz�G��&=`���׸t,;��fɄ-�M���۩<�K�^�#Veggۉ����o��#��u��S�S�B���� 0|�W�#�ۗ���~�&�+*$��ZLj9�:4�8�!G�T�S��7ٟmB&�L
�Ǆ��8���M���RE����}]�R�lW�߮<+>"�>�yX�yd!��X���
?�c�������s�e�R��rX��Q�s��9��3w��)�E&�aQqp?���� �5#omMG4���E+���%�?D��x&0}M�d?�h6G9��
�I��%'2�j$0aHj����W�t�ϓ��0���:!|���Ԕ*Y��g>h5?�̦���Ŧ'
�:Q�εg'�"�_�,0�[�@��\>\v=�,ϑcǅ@�chB��a&X	���O�]>Թ�QK˸*V�c)Z{4�-ځ�?b�m����6���tE�BD$)�_
�hmOMi�H�1���7^�+@��Ƣ���'+yv[���$�_^�&Z���n�ݑ;/B%`�%��}��UZ��ZN��k��k�Є!k�u������Ac�9�z;EÚXD]� �}�͢����Ï����GD>��]<���-f���m(�-�)o��?��t�����C���|�34O}K23^��D�;&b�v���T��E�M�����Nf��D"�K�o�-�;k���F5C^��蠲N�2�^�8�U�H6�f�����y0K���ڰ
/թMG܁�z��&����[���d[����)����.�6Vb���AxG��YKl�W~��wH5 6��h�D�L��jV>=��( ,�z��o�MR�`i�Y�[����ad��j�HS���M2b��[�xg����Y����3)F�t����eN�ZK�%�~ �w3v�eC��?�ʞ��&�\^O؇�x�r�:X��XK��u��a���3������[ʀ �jM��K�q��F+D����|iAQn㡲�ڽw�����ɓ#�1�/Mg�O<�;Ӟ��36�c���#�߻~��_��k�s�y�ʶ7~��L��u�w�T���Tt���s��%:�Q�M=��=���Ԏ�Q�H�9��� �'�\Ȣ���Q�p@���� �_o�H�n�/"b����v��*�5��>�f��S�k�V��y�:�W-�R��_�AY��qxxxZ�(�Q�Ry�������A^�����
G�[����73�3�#���7���N�5!j�z�r�󧟣�\ K�^�eo,ӼsЙ����3R�|j��j> �uW����N�`r�+s�*�Pur���#��*1�h�]��+ a;@ݝ����7�8��h�!d'�E�@\���l���On`��^>��K�42D�z��=T 3���l·">,&�Z����&b����a�#���o��J�ť�d�\J2Uq�f��jL��3-���Xz�Q��2�[��<�C�Y����Σ�*z����ۓJ11~/1�ꌛ�r�Z� Ֆhf��*4e�h�P��Ɓu�/��C�f�B�?��o���Z|� �m��M�^��)�7ɗWuum��~9���˻��֡��vl�<l[��$�S�e�+ü4�z�ś2颕�^l�.� �U�
*C��g�9:��jh��yB_��;(����7�CP��M(s*��;� �5���L`}ZќM��|��[��4�
�����* ����_�i���/�ͯ�ٺ�a��o�~[g�(�dP��Ö��m���6�0���xc��_e�Z���|��ј��C��X�4�FJƄ�:I���S[�\�z�˝�_�����}UqAՇTtF�V�l�AF�;(V���4�uǒWP�b&�&ɡ��c�V�4����{�� m3H�VW��*�ÂR�z���VX��� ��k��׊&=�"�|4r��ׇӏ:���3�$,�N�@���#e�����W��y�s������Ҝ���q�0��<%epz���+�߈]D�\�OqU�X��3��a�QE>�+���ER}�J��9���R��B��G����c0���b|�GqV�z��]�X.�0��8��Z���U�1�o��+�˃�i��ʷ��@�����Y�㖐�o,ٰ�_"����<ǣ���*�M���,��i��	EqQ�H@WH����{X��ƓO����P�U�uum֡�ݝw� *+I��9Ľ/��A���I���i��s�v�G����Ɇ���_y���.�x�9t��\�#BV�|I��R2�������!/�7�j��G����ΠoL���������8�:�%�4 ���LH�۴��SDM,���+5ni�-��8����/(A��5����,f�3ʤ�ʪ�v�����p-��喱Yl�?��X�C�;sV���N������l�] \���&أ {(��s��j�Z�ϴYzݠ���CV�D`.�Ğ��'��8��}������$�c+�F���~�����~סwU�F�w�iC��\>Eq Qד�9+��}Yh%3�/�U��^Y�Pr'�������c��:�;*�\�0n��@�d�'�t���++b}]�?J���[���j��(YԄ���k[�w���E���%H����I~��/�������ͺ숙~�d�﨏��L�d�%6%��/�*d1'u.9�|�aFS�����)��YA����d�? ���>W�)E����t��x�~?ow���#ɳ�VÊa�`��B�������>��6�9$I;������?�뮭�����Le%wq`J�~�d�E�v�-��JN>0>�Y�W�r�[��X�~O����"����l�5#G�83k�{
�Ӣܛf�%L�?q�|����~���)<T�N�J��PG��Ki3�����!�/� �[���D3ؖ#�}HL�3�᛽X�����Q[�n_|��O��!�>�v�9�ilSb�����@��y�-fI�33l�wG�;�j�����s�?6��;�bV1��#���y(ՇRfU+LJ'^"�B��vk������B�	�$x1�uy(j�`����nce�m���a�Cf��l�ڿ���2vӠ��Zm7Z��H_qZ�P���د���3$�v.���.�SU����;�ĐrD$}cٷ&P���y*x�Lw!��rlHL��a�8��>�tM;V��͍��D��W�c'ݙ�<)�>N�jk*���%G�8�4��wR��w	l!���`dR�AW��$ʿ-&��f����2B�������o��.�����_uG���o`YC�M5=��$�z�H�.bS�sC��e��/�Ї�Q��+��+�wD����l�k����'0��C���\!��P�)v�{Һ��u�S���,�>F���}�B�� 륧k�$B +�-E������>�j�A����>Þ��a[~�����ǅ�����]s��~�5�3�UpY�xw�6�	M]o>rh�kV���:w����pu�l���Hxe"oؗe1%��P'U~��4� �
��g*�&���c��3�b%`O3��'��y~��TOl5{3���wm�s񀟯$d��*���6��*��Dx@UW�*�P}�5<�)[��1����Ow��u�]�LH8ӝ��!j�%�_��ܗ�2�`՝���tԀiv]�C6%d�K�Շ�H��zt�w���Q����7�e^�.^[\d�пEZ5�<j�����IV)�ʊ�����$�<D�-��_lB��/3{��"�0��bp"ry2+��A'���K\� �jNy��:�H+:��蔳EQ�[���T��q�n1s��rx3�\��W���o���R3`��^�~r�O��5�j�H���Wj��w_����?t{0Jh�A��+Xh��L��`1}j	��5z���'�A���#�c�d*� 'A�\�f���#b���JKP���Z��9�վ���'Z�^�/.�98�r^md������2�x�.�n�φ�������YG�G�������'�)@9�����/�@)洆�D�)*�CB<��O�d��H���	�5��ʀR'|��uZ�%^q�W��N�X��n�ⅨXt/Cg�bݢVp�[Y^t�+m�A U����1MF��&O�3��-R��Ӽt7����d�4��aZ]���U�Ȧ�B�c���{�Veo�a�H��J\ȣ����oRk��s%e�[qi�%|'�;+�3_rX�
"vGNW���|��7&%���ߤ��k=11����m��:#�������?ox�+8�/}�c�}ߒ�튉����\�*��A힇چ�s�033HW�?�%F�UZ�k��R2�t����CC�({e������e	 �}�s�Gwj�S�f<�ƭ�$~��O��]��J���B�"�ɷW�O�ϮAM��i"�sv���"�yS,��=r��s,�L{�5,*� �p�  �L^8�ԓ���,B����*_�7�4��/�3����42M|���8�8'�+9�6�%�λ�/�z�k`�7���]��J;|�S�5���A�m���������u��iR��,P�&��zR*�%"���B�kfjI[����c�'����B���<A�T�°��${ǩ#s��ܞG���3�U����1w�L�x�\��B5"�mV/G�]^�z�2����o��|�g�����si����?��z^{�B�%z��]5�+��/�iXZ�T4H&�ht���ڣ |�Y��x���,���0PG;���0r��i��2�^��l��x�Jv+�O��N)����T���<��FP`��%�o�!��&���Am��ky�%�߻l+�8H�l�
�/��Uz@c,�ư5!�8���52ɣ�����UEX��ӷ9�˭�,��M p~�4i+tకU�-]#�l)�GYQG7���Uo�>}Q 5��M9�B<�J�0�d�w�8��Ȩp4�:`x�:��j#���^�A�5��Zxe�IďjM��s�ƹ�=����x�1C���"j��dk�oӆ�j��S�������^����l?��-5B�yW����KG�5)R��r�`��XxAԜ���	�����wrN? ��YI2�����L3[�r6��V�u�?^��A�a-���R)i{2pS���f���~D�~%���
��(?V�s���wS+�����_vU���c���T.)W�q��`
)��oը���ϯA��s|�Dt
AU����%@E�J�,���U�^��39�t�HT����v��<��<؝>TD��-輄�m}��Lu=+�]�l��T�
�ɡL$�u)#EZ֎*&a ��� ���?��&�'��X���D���g�j�%��o��	_%J����D667� �� �];�=��ڜ
����/���E��VÞ�y��i���~��	�u��MлFz����W�4O�.O���eӬJ���9��b{�/hxfh��)����wp =s��c��Q���n�v�a'��)!L!����ϗ�,���Pwi��6_�dD�)�5 ?����p�X��b�R��|���!q3`o�ޅ����� ��]P������ya�X�p ������SI����u)|�c_�(�7�#������O���
��zz��(���P5(�X1�.�bU$¡'T�-�;�FE2ь�NM�$���>�UV�w"��[<s}���d�=��rW����޽�Ks��V��D��{ܕ{7�h" �ń���{%���^�r�i��>���0�Hr�JM�(�[4�\<��'�-=���=�&��h��l��aLs"���?�k��~1 z����m�*l�a1���?�醙=���n�N[�k�Y�e�"�x�U2~���O������A,��G���x;��nU�����Z��˝�峒��)�e%�l1Zܛ�Ȁ���i~7I�T�2�z7"�-� ���C�
��_蕼_�����0hU��jv�� �������g�t�Ǥ#P��󿷋(dǌ�\��rU_�P�J:�qD����'�<��H�U���%�]�TUN�`='�T� �=��0�
�K���c��6e��Q��'�N�+�J�!�c~����/�1�rd،p^���"��&�i��pcƐ�ꧡ���K􈾟=��{�@�`�Z���N��,x��������p��%������̻wr��ܹZQ����� �f��aU�K��jcL3@�̟, �U0��L�k���>�YĆgTH�w����*K�p�n�=�4$E��P�㷺l[UxFtlp 8WA���Y��-��g<e��yNd����$k��Y�ӈ𻆉�(��͡|�����v���"��ѽf������
���'ݖ[�'�I/�oз��wV�s�0��u�k�ul=Z�r�u̒���	�K�O������{�z������m޻�,���j^/���3�<�}�Y�OC�ugm�A*D3�8����q�c*kz�Я��V��r���lR�{�k���/�sa�+6�t��8ӎ���ƔR=o���o�)�0W'��q�!��<�ז�-�8�,�����;�|��P�l�g��K�❱�1]h�4ԻP�yK����>�[��/3�������Mw��I�l�D�>s������mp�޳�59������r]5uuKGG�TU���|>T�U2��ꢟ>�Ud�2Φ�����Z��l�
=�K��T�4�Э�p���x8T�w�b�&���D�\��4#B]8�Ӧ%��y�A�s5.i�n&�>mU'���5��j���'ٓ>[���j��C�{\�d���a�����#��N^AW�nvv�:��Ƥ�ώp�Ʉ�s�V\�櫛�\ѹ�w�[���_s;���Ͷ�����!��N��W�P��eb H��R�K�dd�.�T�ȕ6�Ȗjk���ՙr]z���;u��r�	�&`6��s���ɔ+Gz9?�oc���L�h6��5�W�iu���1�t�Q�:2��'��:s��>��a���r+��9�OBU�n�t��m�,����9[^.�5X��e"I���)5�;��[s=b�g�\�M��L`'��ʚ�bᜂ�~�c'-��Q#M���Cb��el���?G-y�a�E��������'^����QQv�ޤtJ���t# ) � !�"%� Ҩt
HH#��J#��H3C����u�\�,������>g����~�����w��qț����Q;����kO����[�$oo�������K���"�|K�= �$}�52%�nw���;����eec���UϜ�0�;���0�7۵�����A�����,��MT��~��"MJ�Ŵ�ʮ���S7Ѯ��9�˲)Ͽ�l"���#�:����aò�sM��fb�����ô����Pl>~��S8���63H���	������6/�:��S{v�EJZ�.o,Yf��i�#`'��|�QG$J�J�'Xc��\��d5��#���) ��K����Ff>��}� �Jz�7�X3�Gk9[�"_س�E>f��Ń����]f��𴴴\dZ�Vs܏���n>~l��,��a� ���ii���%��@��̖Z���xD�R����*"f�r�b}�-R�8��}��Q�(s�!9�)�۽��ז�8
�Ƣ��.�E��A�������>�2-H`-G�tF��($���w�|Q�tGw��+a�S޳�P˭NP������hL���Ԣ�� ��Ym�Qm4�	&))��������e�qV������#���^���с�Ч �gnVu7��ƫv�O:T)c�Q�n@,��\�fJ�H=<<$A�ÙOC�i���J���g�F���fJ�ah����u&~��x%&_���}d������s�ǣ��e���n�<Z�C�]�<��c�rE��褁��V̧�Q���pU�i��3ㅯ�$��4t�G��� /��uyN��eL�f���6"�OMuup�f�c�K��(d��<OcZ�Dٿt�44;�ҠW�/)�̄3o��T����T�^W��2q���Z�tKv��6�՗s��f}b�@i~pr�����rfaNk�]�f ��2j7ˢ�C|n�+�J%�/�4�e"�+4��-�%Pn�ʆ��7���^;T�jO�trf!_7��q��I�s`�m���ULrQ���|j�Z?F�+�0�-����+��u���[�'�9���?g�m`X�O~���z�9�w����܁9]�����s�*Sh��U���|�s�D6�)1��b�[+��>Z��b7��k5����X�9��o��k�eh���0��Pk�?��D&ઑ�$��ۡ�!�S�mmquuO<�lV��D"�ūm��UU�Oͧ� |Y�#��o�t]�F�ܛ����L���_ m����o��j1F<���+yLo��Jj�'h�_��ԧ����3z��7H�$�F?�]����^<�D=+s��'l��w��(¶S ��"��5��ȡOG$���x�@ȯ`�����>�%_��)O��c��4k�D���I�(U>�
잕�;���X��,�N˿�Z�)&��cҍY?�.P�g+���Cͻ���d����_SO/|��n�c?�tuu��^����>h6���Ԅ��ޡ��u>�WCS3��sn�=�A�Y�Q�^�-^�3vK�����@�Ufʂil�3;�����9�^V�:�N��B�}8��YT>i'��怲��A�!E�x�-&F2�f02�e�/x�
<�7��c�#���u�1�����;���>�Pbt=� �� zSXD�
�1�/��X����67�.\������nF��(��<��HWF��]��ߠ{�3a��@� 􀞞��x�bjj���9�/�y��@�nY�g�St�C�`�@jNN_��4:gL��莎�]W�*L�ြħ_>�)��`~�jÇx�9�����_S��wV�J��d�AZ7��ٞ�*���~���9��b��Kk<���q��M;��(�b��%4Z+�mt��ay�ƶ�gE�������5�N<#r*@�T��.�\1*hZ�L��UiZ>�DYZ.E�l� nĽ��M[�oib�e�ep�,�%�7��[�����M���d|q��_  <<L�-�Z��@7&��� +,Je��g367ﻸ��%�>n����Y�' iMZ|(6GrPp��GF�M"����t��]��h�g����HI���h���:Z#hF����A�G,hAY��/ "�(����f���lŵ�g����׋1�x�,��p^�%�E" ޘ{h_V�;П~k��SnI�F�O��A桄 q�v�n�+8�nL���|�飈�>��w�]u虁�3������66��L�y˞݀&605���q�����z=�1l�A>B��T��1]a�Un��z��O��F�-���#�S6Dx�����W*OВ�2YŃuٖ!b3V5*;�H�}��X?��4�����~�F�ֺ�8d�����}�S��c�ZksZ���<'ǳ.j�l'��˝�J�S���������>�r{��c������^*��r�g��ֺO�6���}"]A���3O���D�f�̓�`�吻^+}�;Nd#:Q!~�h^mF�o{J�k`h�17��I�#]c�/}�X�G)����)��?��]Ox*���x�+�C)��{{{��2�T�"�U�b�S��`�Xꅗ��\̧�;MJ�j�=�o�}>��J�1�_��{�>��*�<pd�,�e���a叝��|��$~U˿���� 	~�����b������`��қpo��^�B��%T��`�=�!"��Oaܟ%��9���Qr�|ի���ᡈ��>�7��m %hii���-'-����X��ֲ$i��o�f�rC�u�K���Zo,}�����|c��t���� ��F��CEQ�FɽI���ū����l��?�y�Z;-CstAA��ј��7Y�Zw�Ozo@��ˣ��C�J�ls~N�ƚ55�2��~��C�rys����;z���@�O�(�ڐ�� r���đ�;�E�9��Z��&i�o��Cȿ������#\gD��a���������r���wAe�k?sO�M���F���1A�t����,�JMH���Nhe���/%��Á�����ttt��<�4n'V�����Gypx8o�é�M��+�N\�z�<6C�J{,����N�A�rV�
�ɓ7y7�Ƙ8	>��*��x/SD����Ҩ�9����$Zܺ���AOi�$����=`�Vf̀Q&E��:7%H^#s���� (X���M�8Qա�;�ڢ����v;��/N����^�&f  �tG����4r�t�����f`b�`j��'���P<����s��t��7s�Е��K�r�I��vO��oZF�LUܲ�c����l$^��_nk�9l�nT,py�:�ȥ{ѝ0����\+ڨ�
p�n�~|i ��hG�e��Q��y�=��WeQ�L���g���۳?~J��}�nnL)��w]�����%�������K��P�w~/�Q�E�cZ�R5��+����^6�{�ō���~h�������$Wpct����Oԛ�����f �	O�1ȀO���� ����INIA� �D7����(n�ۘ�r`�%������H�p��Wfw����i3�+i[�7V8K���F��_�џr����h=�v���	t�l	8�ep�K��COXxE�O�G��m�;a=�@2��F���uV% �~�[��%ߗ>���c=�`VL�2���)���:��R@�A���%�γI��P�/�^>MA�#����m�*����p�V/�}ח(�?�9ܢ�����H��@�q�L)/B��cJ��0t至�}��S���w�s��v�PN��p�q�*X���=t�2�8K��l�Y��H��|���^�^D=�gߓ�����[w�ۥ:��";e���Z�k��j���K��5�z�T�f���N2~gBcsJj]�Oh� T)M�����_pnb\���-ݭ��L��y9�_̅DD��RgȖ��(U�I��9��?�)#7�aNh�$���Q'j)p����Kv{7���R4�E0�[h��<?����:�Y	�u=���voڃ�`�E��������^��MlΣ�~�]��}BV����"��~#�I��%�U��6E�#�s;�q52ɳ���yG��`E�N�����I3.��Rh��8����ӿ��j�u�B���G�<[˷,�z�<���b�;ńz�6����ɴ��2f�徴�ѐ����L�&	���M�s�g(�����bk4��ň�����m����h9aǉ`T��bum^�*���XX�2jE��C�,j�S}8x�z��NAꣃ��W+�?:ۦCͱcIb[M[D[�����&5��j^����|�Y����7���	����򙥚�������b����b+���?���i�d�>��������>\����*��4����1��/ƃ��]s����\�1�����O� 	neoO@DDtv
sAF�_a���S���ښ߲�����Kk ���םD���_O�]��kQcHB�������o��\�>�]�uchb�6v9�r�=���`gh;lv!�Ȟ�i���������.�M�,!M��j$�"��;��l��j��^m�r�v��W�/뙮�����S<i�@���O:9�ϾȪ���Y��6?�9Io��u<ʬ4;���<��I����� �c'��ߗ%���o�<�n�71�ۥ53%���A��pX���ry��xԫ�]���4	{,]W���'�ª6�L��ʼ�
�^�����5���0�@]�87���Ah�ǁHP��5���M:���y�(�v�m(_�.��I-���gE��6�2���w����MЋ��vpg�>4)}����i�MK�S��fg�ox�+��kvN���>�D�ܙ���E��:�����3�U����w|p�S�l�8�7,��\��)�uF�?)DHOQ��N��((���oֱ !��	� ��l�To*���$�ഽ��v��7��-���=Q��Z1�����P��}ޞ���$�Dm�ry���8n�\�Ϣ?��%���{�������Sy��"��*��Ȍ9l�%>=�t�<c ���\ox��:�������S�r+ƪ�>,�zB���g�.G�ss}yvs��4����O�a�ێ6l������4�z�T��>48��oӢ/�옂�`�~��<yA���`�mgC5�;! %!	h����X�G���}�� &G������������e.6lm(-��dI�������^�0��c����uO����tbYe%��.�ٿY�u�N JK���f{d&��!ٹ?A�Tvd{X�_f�M�������/��6��cjhW�||#�)#���`o��-����V3"�55��)���hU�Ԩ�fF�cnݐ�MG�Ю����V�ǩ���?>�=�yJ���5Ɔ.dd@P'Mz�#/3�s�;�������W���=��3��%	b3QOڭOV|��4�^dț�i�"�q�,�������Ht�1Q�y^�M@]ԏ�����M�IK�E���=�M'<�<�	�~Zi����1�gs�L*��� B~ڍ�d���#QMMM��.����=neee��b�;�+�-��5���OK��Ùە
��W����hB�>CJ�wW��
���-�t3]�	������Q�zf���{LWm���ee��}t��}p��'9^�����@�W���N~��g(Dk�j�]�����]��W-7�,��⻊=Z<�����떖������E~�������#������c�LXO���� 0us����=�~KUU���5`7�I�T�rc����;��y��&���m��w������R ���Xy�G#�(��ió4�A���c���x�f1��Q�tKU�^䞴IVM�7� әL���1�K��ǺW�Y=����wa��G�e�I�ʪ�Q�sjm�vn��:uD����I�O1qh�p30�Y\��)C�! LЮ����x����g����	�o1���n9���Y��� ZP���g����Scs(x����"��-&��-�7�u6�����k�h���G�1�ЈH�,��!����s$_}q�}w�Ҕ*?�����^�zD��+J�������@���O���ݲ;�+}(��\�����!~��!���zB�k�Jp�S�o�L���Qd�U���Z�*���=�S��f����L@�W��4�w�_��-�`�����j��Òq�h-�Ǉ�u3,�{Ⱦ�w��r��q����޾I�AO!�M�Jr�%C�D�?���_�-��� ;<�7��%���NH��=]N�����8x���c���ؤ?fXnoq������Qߚ��gU���L5N��7��\����6A'�Qu��x���9�w��F0]��oZ���:Z�̇�U�D
�T�o�(��w[�gp�@��ΰ��9҇
���#���.�'4w�s2e����=2b�-�^S:Y'��/�Jg��7l.�cuɞ�kP
U���s��N[~�:֏�}������1�T�y$�o���_�l[��f�KZ��ze�6�[	~�Sc;R�4h���@�����L�o�R�p��/�`����eHN��;�ݐ�C<w/eCC�ik��Y.�M�6��,�!�Ŋu�J��ٶ؟���G������~H\t*�_Q���ґ��n�R>��!�h�Od�W����^�\��| 9y'N�����F�Zb��U`�i�(�b�Φ�T�������_��my���&|P`�M�P�K�*v善�yź�er��&��9���}`��z�?�!�XhqĶQ�fc ��Лr=<+��U��
����Ϲ��N-�M�+��-�y��/��}�����ѫi���5It7�(' 
г́W�uF��U�q����#�,��L[����e�%���NP�'֖�.���FKԷ�͋2E��O^���z���XI���T���GL΍�&^���yէ/,A�z����ux�eAv�$����{Ƨ���"�~=)ƱE$�/�� ��|�(2&oo�������y~o$[V�%��2�%��A����[DOI�@��8����j�H� !��C�a$Kn-r��-�t`�.Y+�_��� ��������ȘC�;Nv%@!�o(ۯ�11DEE}.��ai���R7oeV���њ��Y�ou���ߵ�v�����Ԇ����o��-����k�5�Z�F��#�����g�[P��{ň5�u��� �v#Ka��L%������њ������r�痊v�	B�.6h
�WK�Q�`�9�-����8�D	6�|���@���_mH�w��Q��2����ƈ����ux��e�E1���K6 A7+7�skq�f�����)o�._^�1ږb�l�4����AK�z�`���0�rn1Q���r��)J=Օ��l=KM��&m��!��b������	$�.I���QXT�1���w�i���V�j��x��B��rR*�'z.��H�9��U@�`lQՐ!8wKWՔ�$cN�+��'�uƨa��ɝ����m�ݚگ�.H@Į}Ք똚�Cgv��C�㱗g[����f���^�1_S�^{]���dw��5W��_��)���#������[��xv��T�-&7VT�Qlz4�]f�vA�J��{Ԯ�G݀];��<q�u3@����!���U����:Me}����C�B�l�����J�!ᛂl����G!*�(�fe#*��{~��U�(�����Ct����� �HH�k��"a�B33�������0��m���ɼ��Cd�gJ:<�kP[n�����.�!e�y���3�!� �}tg�8F����%*��b�����7�zfO�]�cM�>�-���ϩ:-8a���~���CԦn�1�f�*��z������p'?�ۀ�Ҡ���oNѷ2 >�)�zoQ�;�ēT2"J����|���\^b`��Yf��J����7�5:r������*+��+�F�R�t�_a߬0�`��&��|�!1�3���!�,��n����G�o���V���\�{\`hi�k�q�K�!Ѫ����j��:"j3�BT����cv^�.8�H�ǌ������,���$j���[[���������|<r����Cd��ZE�u뽚�`��/���}'�)�a>��s��v�����O���ؖ���U��ꎠ��z����N����b��_���J��"�J�W����m�)�X~��z��a1,��[|Z��-Z~�P�̿9Y��ߪ�Ř���P]�R��������X�3iV���{3���āWk������o�))uW�X��ࠗDd$:꼠��O̬�u=<U׉u�d��Meϛ�&�H��T�2Ƞ� _�ۉ8�MU��*���#�����M�E>��Zܶ����I�5���G����E"�3��c�]��iJ2�o���2?ӟ�\E��ߦ�q1O�x?Auv=�q�U�dUעd�G��\�r��/����M���5i^9^�ݟ��Q�̖ `mq{s��E�o<d��3ݑ����f~H�� �I�����*�sw���9��$�O�x?Ӛ�;�S���pU0�J�q��j����O@rm�$�J�8/m8�����Q�i�|G;#�L���r�� F&����Tw�Ӝ[|����}��lH��
6'k�\�p9ܷ��U� ��O'��c$N��'��Qc=5�(txS%�A�X�E-��`.}Ukn��-���ڪ�)r�~u��C����ׁ�����ؿ�b��x���>-�����KA�����q��.�+�����)��U1��Sm�q)��;�����4;�\��d�a%�Z�O�hꊒ�֗�Lx8(*�qkQ�R�2aΙ�>n��I��ק���*�r��S�����+Vt�b��� ,0�R�s��b��ѱ;3i���+�'�]B���� �F����?�M�W�E!�~������֜�8���,8+=X�P���L����&=M�j�^�
c��I��d�t�[C<w�H��g�僕��[�z�����x����ߋ�����HI���^�v�7To��#\%������SD>�1�5�hee���*w�Cs������?����d:�ު�W%6M��g~��ڢ޹��9�<�8������W�j^\��)8���G+X�����H"��ܶy��B-��rEz�WL�	�,/6��9�R�rM�_��� X�/�^�:n�j����	��7.j:W��w��`~��f��'��[-��������?���������(+4e�8mgV�~GCm~O+�.T�w���a~�%O���G���ˬ�Rߪ�N����3��̇��z����dy��&�k����I��FF��IŜ�)S����)����.ϵQ0����`��f�ă�����?m�}�S�uj"i݋�����؟`"�'D�5�1�$��<:�^�( E����t�d�����b��b�5f��Mt�������t(�P�=X��)���	6�����T�=S�����إ&�
),|lx}�xs�[m�C8����3���C
�Vf��jU�M��[���`�sm��r��b7�*�>�_�EY^���w�7�nj|�Nl{X���N��i!�ǟ�����s��@Q��F�[�f�`�e��b'��L�P',�LS�R#��)�"�����]{V!d� !���_-��+:cF���u���e:��Ԝ�ِB��s��@���'�f�^��J��ճ8?\G��/�/ ޛ���I)�OX������N�����^x�-��G��(��O��@�X�����ß���f-r�o�`�'��<�+����8���W��Y0���u0WT��%��ή8�f�4>WR�������ä,Kه3�ey��F?&��(�JwB�I<g�Ti#_=��Rt�Tx��v$�'�Q��	&��������P]h�����P=��~���?N��I}�X��5̻���J�f�V,r�l�1B��yx,	-$ ��'d��N�$�y�/n���3l�	�M_�M���,�ݼ�B1�W��'����D�.���p���T�C���>���J!�C�v���S��(�Ɍ��7��w�2��u�5&��Z�!?T	���;Bg� A ����[�(?i��Ӣ)����Z����s�:�	h��0�c��~��&���zc�<ztn�C<zi�����c��h*��3�'���/:x���T؅D'�F��Oʹ���E��^E�,N��*=�F��p��k���^�.2�݁�V³(��oS�ܶ���A1!wi����1�=c��x�j�:�C�Z��x�^��������9a=x����A���X��^7���#g
����0=�	�H^Ϲ���ִ�SN�M"�����G3*�Ot�L���E���!�x��������S�z*�A�bl@��a�-gb(Ѭ8�Lp��ޠi#=��B����_Qe�3���#��,.�`TŃCD:�!�|��(��o3K�W�>\}+���K�G��+���_���B�tO�Y[���������B�Z.�p��o�yƂ�M�����WxC��"���xB�49��W�W��<	mEn�����c9=<�u
bQ�����s󌸼�v��n�%�*���E@�����̋�D���co[
pCX,��=�����=#k@'zeWT�!p�� ��܎3//�y1.��&��Yl��m�Q���oi����ʳ���߰�UN�#����bhi>���_�V�f_���Y�U�t]� e�2�9Li��9P@`�A5V�Y7��Q�����O��W��Ab >)�h{�8|^�g����Q6ч��n��f�lY�Y��IIP����d(�fe��P����W1��3/��y��o��rx���apOQF�{�D�ë̇���Do�����N62\���I����g�kS��ëv^�*3n /T[�1��%�D<IUQ�D<�9��!م�Te{�%�CĽ	`�o����hR(}�B�����&�
���0q`b�×�"��ԃ.����#
�?��/�ݨ4.��"o�B�4���^���2�:�Y�1�|խ�6�B�/�lE�˸�┲|�~D���{�Q� �(����lO�ݙZ���Ns�I���یc����*�~N"�z�=�sj\O6�"���=��l�9����T������s�w�o`aV������ �R9cD�a]��)�n��y�L"d�����&_:�8���h�N@{���Yp�f��ч�l��(�Z6��'��3�:�N���(�Zh�K���A�t�j	 �)edḽJ�X�(���16?�&j�
�n����Ҋf�<.������N]~�\�u�##�`q��61J�܈.��I:|VY�-t�!��c&R/$Ȁ�y���:�'-�<������B�XxF��$^���_,]]�?)�W�w� �e|�l�xӃ���}��	�I��Um4�U�LC����߄�H
��S��D�;�u	ݫ����@:g��[KII���� ������`	���ѭ�����_��U1F��J�0@��)狰��|�E�:e	��Df��v�����������E���]�&�e�mMCj����d]�"�.=�mᘘ ����N-1�YHԛ������vG��w��|�SE]os97���z}m����sP(��f����yU��䫲���>7�H��Y,��6K�6����V�����u\Fi韏��4h2F���C_y��gzD�k��K(R6j9@2�/�����}�A���͵�%����g��XIrb$i��{���u�;9�b�����{%�%\�"���1Z�M�ۊ���� 	��� b�XQ\�Q�/��͐�[��j�H��U_<�e*�����+++�\گ��]c��A��!:�������쏄���O����-�E�bh�.4�8�W�>��m��=���'�����c��L]}�|�_�"�<o�/�8��J5���&",�H����:�E��@A�'tP�	Ff�}����+��J O���p�[���4/q���	]7�3aq9��"T�g%��d�9�_���q��R@�چ���^t��ϸ��z���K��i"��l��q���%�8B�yYZ�C0��������B�{���Q�O����bp�(�p=�u ?�Xd b!fIf0=H"׾�aW� ����љ�=v]�PW���ʤ��� ����$}�;,��<�ʕ.���*'	�XL	�T�*���|�T2f�T;�����ڂ:f��Av�N#��s��_@[�M�m��<���*8Pox'�U�4}����O^=���Y�{��}́)�}��Q0�vƓ��4�Io9K������<�"Zm�#kV@
�?y���矼�AT<J}˭wjH5�ҙ�-����ᒬ�8��ae�ǣ�B]�ʓ��R��K��Uy|�����"D6�fsW���g��j����%�?C4V��P�&��ԥ�Q:�O}�@G��}%�K�m��b~x3�nl7���MqG��i��H"H;s�"Jͯ	я��F?�O>l.��<^~28�]���"K��y<2�t�к?\t���Gz��mY�ٚ��R����/+�s� ���n���!1�!�̋�}�5��D��}�o�4Xib�f����)��B��*�� b�$�
2<�3�_�Nt�d5u�e�����3���="��sOW-w�%ۅ�g�s�(�mn�tSw���������x�i�J99iD�����-t�~s�95��I��:\pRs��XK:�w�T��2��6lyJ�vt��K/�
���+�/�����/�|Nb�o|�'wO?d���"�C�=W_Ա�jpt�r��[7��Di�����eaP	ٴ�T�V���2�jD�??�i�LU��Ej����?�����t���Q}�We����%��@ �xcw8	����X�\dJ(J�cs�����h~,-�r���r\�~ɍB�'FK`�gK�A������T�h��`��-'X��(���\�
�n!�)��餪�V�QV0x׭����R(}u+��������o�wR�_TD$���FIw-�0����-�«��W�9p�Y����ӉZ�c� hP�����5ml��T�ת��v��p,��z��l��&djJ���]Ĥ�yMMtCCC��'�o9Ҹ#-Y�8�����3��)�k%�lm�B��n���))5� v~�Wݖ;�0Z��OʉE9}^a��䎚*|�Ӟ���z\Cq�N?�X���Ċ��y�+�Ԓ�hP1)���o}�b���h�m�<�z�Ѽ�F"���O��|�q���&:�m��#��o������]*�ݒdz�O>P��魂Vg�μ�w}�~\j��d���:v�s͕ţ��H�A�*c��?Y	HՁo1�sBx�^���c����M�x�������:�"BBA�x�,L�׭���Y�'�����r5�B�Q����8w�_}�r���́_u���z�mN̥�{D�ſȟi��$=e���I@v!��ܮ��dN&ޢ՜�fȪ'����m�\�
�Tl���nu�?�tY%p�g4��0}~����� �R��[*ܦ�\&w��7a�����e�GO�f�c�48��+�>��?0�Ls�*aـ��u�,��+ޛ6�Y�4���d��7p%���¨~�������	�zKr0M�ރ��]K��CRF)�R�
����?��4�O�o�9������o�n��n ��!�9D�+4��4�)��G#�a:�I���	�r�H"��S|=�@z=��h}cv.R�؇r�0�1��I�k������0��M��*�������������)�M��J�er#����bI�&���#�ϋS����K�b+�{Q#_ԫ��\w9|����w�0�V�d�wުW��@�j]0��7������&��oV�xk�4�u����_�I%h�_"Y��0w���~�m��b!�K��1C��+��e`�3���E����|�	��5��EP�B�ʷ�b�`v�������H"�H2�p�p!>�S���~��z[��X�©ߊ7حd�W]Be���u�7�T#�Xs��X#��
i�Vc%��a�\�X�Vթp������?���Tx־�P�?i� 9��9�'�����/�
����ޥa)�G!,ϒmF�P?���$�,]@�y�+�eQ󡽽/0����-�<�l~��g���57�q�s���={hm�}�`}Iz�q��#4"�K�������T��0��u����/ة�}~&�V��N9qs\��oq~��~D�X�.Ǯ���A�kĒ�*������&�V�;�:#�cTr4���܍���ɧp{/����e�УR�Z��h\����7k|0�ü�A�H+k�z���S��ܦjbX�S�KK�����X}\���|.�T?=M����N��o a��@�7�&''Yi�}O=6�Qf#]>�t0V|,��+�y��>�������18!?��Nӵ���d��n���ɮ����2�Gy1��۝�d�t�m��}���s0+���v�/A��}B�mx��JZV��Jr��$i�W�9�u�,��K\��$�L4���bD�Q�,}�Y���E��;��¬l���Ȓ�I����NLFc2���c~g�B��ɿuuu�0�l�{����_L��͆x;~T.��NON��lc	n�*<����\��v��{�G�[��<Wko�����w�`������Eد<l.:��GjO��J����o5q!�m��;~V�;��/�ޤM��G8��#qv�3�<,KE�ȰC&����?Yu|?D�'#R�����Wq#�c!�� ��f��T�a0�W�0�$�)vf9�:ڕQ��6�� p�+���@�&7�5?O���H#Z��WGe��|���؅�lC�n^__ch3��1b�/�.!PEO�\�l�ͷ5��E+o��tf·�"6��P��|��5���3��}�:Z�>uͱ?�|s�:���|���E���)fg�<��W_�z�L���	��'�,�	Z�sף��.�`߻�#"ʈ��!���0�~.m�9�ß!y�c�^m����~Չ�xO�=Q�Z銨���r:瘍�
`4�ߥ�x��1z�����H�xT�l�V��w�k���ZO!akgf�A_է.՛\��'e�B�9^8��b�l:���U����M]�Bm�p��*����^�
e)�o�ȹo&�~
Wj�g�K�h��[�z����aP��Q�@m_��"͜��I�fi��w��	z��t\ ��#q�y��)��+"�x�V|*@�;��~	>�iY%�[%����ͩ�7�NՏ�k�3��hk�;U�5�%�5dv����N�b�737'���`U�wed�m�>��e�m��rs���ZT�'�v��n����Z�%�M���u����c���u��&�z�,�:6�.a��8�nاD�JL-e�uև���/¹+����̷�r��h�غ���C�j	=�Nt��]�ga�ں�v\�Y���.�骎C�GՂ��3q-����G%lI��S�
Y�4�ۧ;�&%�Ƣ\5�I�.���<З\�ڣ� D���ZO��� FD�iN#�"_5͘_�$u���(����0���\T�G�lX�+�p�/Ow�Yņ��s\��"��|�G�/���Y�"x*����j�>|���Ŏ�@�Ȃq��I� �W�o@�������+�~w�� �i�7�%7�A������"�]ވfM��\�>�3�Ưg����ZIz�J{�Rأ��g|�4�UQ!���Vz�2n0�)WT���������P����/�ƃN"�D*I�!���DX�����m%��eX��Z��� ͻ�ܓ%s�%�u��d�u����|��!��aј5�jF���}�E��H�U��^5���i��UY������%%�L����P������'�x��8�� Ɖ��ts���1}�'T�E���Y|���͌\#��I]ގS ����g����E��-�� [u��ۈVl ��}7NN��1|�'���,�}I4L$j�J�����>mM���ʋ�����B'�T�ah����`�$���_���^o4#/�g׀#�~�A"�n�~,1�2r}"`m��fŒ:|�
Zb9�>_85�+S(���#\��0퍝`�pVT��%�w��
��)H�H�w���ZT����Z�Ԣ�]���sV��yGϠ�������"cX�%�SEf<��ۈ�M���ܟ1���|}�]�B��Ƿ��>��}HKf�@�cNW�o����E�������#�ǆe�΄�*�b���^δ�% a费��:
=ܿ Vd�����(��h��H�qY��nYW�� ���L6��P�I���9q@~bs-!xm���*�e�Ͳ���~z�����7%�ۛ���o?�6��=�o5��2�0���O�>�|�� 2�b��1u���W��w�m~����LC�?���Q)+��r��|���\�f v�$����������>��֍9�6�v2#�?�sv�-�l�ڭ����`�7���|Id3I������z�kGߗ��]��7����G���Y��K8�#ސ� �@Q��y�	S#{p�O^>�!$��r��\<�I �U�������Q� ��T��1�r�̀���f��,,*)�	D��۷yVU^������C�
�� ���������ڹ���2}�c�����V��	y�W��k�&��4���j'�x��ဤ�r�m��">�; �-t.h���c�#G����; �*���Wb��ϊ*�c��?��#��G�u,/`>-H�1O:
�(�9��(E4,~e%�h��z���X��B��l���%�#,��+�Jņ�f���8�� ��ԩVV5��
ִ�V��p���_�2�\Q�ٸ��Q�=�򱺥z+ ����f:�)p�����|�eTUa6Lw�$�i�n�C$�Cww
�ҍ�HHw�R���Cá}��y�o����u����{f�k�����e��u��y�(��<��d�X��Np�[�E��T�d	����?��{����dƮR�q��S�\`@4�|m_��ל����=��6�S�'ϰ<S
-��h�<:2-�%�>��Yu��?Q�������qw�i���q��_ՙ�S1�j�e^���%Ӻѷ�D��9M.�P����}��ul��FX�\�����GGO�V��,̟|�HS�ϡ*�Z�2tL�<��'�}���_�����5T$��E����'��[n���i_�o��9�h��<�k�6�3<��6U�%5O<¨[V��s &�<�`/\
�i�b��� `��J�߆�K��$X����y�fo��7ƿ/���n6Zs4�3�6b���Z�Y�+6�Ǵ\�C겋���umC��0Ye
�镯9t���я�tg���k���|:��]]��JA�t�LYbf��n�����W�㓓h^y_�����BqN7�*7�0ާ7V�X���V��T0{:����a���	�D����dm�wc��%�7�U��їgU�	�
��p^�~<%b��7Kx�x��_'���{��U�)�X3M./��x]��ml��W~�՞�[e'<焾��e�dB|�|�����*1 &x<%$�]	)���|ݴ�AZN���t��)����?Z 5�����묢��8��0�DfX�!���kV	��SQN���A<3��"8��5L5�-1�|�b�^Hw�,e��3�l�c �q9'RNx'�
u���X����{Eϰ�J�a�h����.�ϔc��EVJ?uCGiIJܘ2���3Ѷs�ul���M���%����\�=B~U�� ��@V��B�wM� �P|ن�����&hy??�� e,Ff�.�u�<W�ܦ/OR:bY���xqY��3|�o���5��b��d��'��M�rmP�d��>M&@-Ԑ�I�G�|w����~p�YKpӄO,|g5��TA"A��y|y�!L���k�f<�.�͗y���gz�w�����n����.K
�j�n�9�kf�7r�Q$����C�O��φ<�(�3C!f0�헺L�2��R��}ۓ�o>�0˜d��֗H,�� ,��?!PYE5$�3������js�6�ߔ0v��~<��Ҵ/��r������i�1DU��T�Ř�#�zBB�F�o��gRBn������ƽJ�Ӛ>�'9��Fq�'�ѴC�˼���ׅ*�>�!����O�+2&Î'��<�ܤ(>{���r�V��,�q��"�>��Ņ��`[�D��7!���ϓ֬�F��/)�����l?��g�}N��v�K���]eP]��GP�q�~ܶ�I���M�X�c�6�Rŏ�(����Ē�����)q'�Ii��X��ؓh	��D��W���~�F{w���W2?䙂vĻ���z�Z�������V0�!��C��*�u���J����za3��}�����N\��&'�����*|6)��<i�V�2�"�bA�&�?8�� �BW���~lm�+�\6��o2��V���1�<����/�o~繯��|�+��,����R��g���h�	L�\7����8�s�?o7���|��� �+�`��JZ����.�Cm>��/���kI>�n�߳�7�������Dp4�/�^h٠�� .Aclhjv*u�K0N(A?�5��2�u����Ӝ��J�zfJ�vhZ���f�iZ��nyC}z�����^��Pf-�w����1���m��b0j�K��������t���v��{ގe��w�	7��4Ьȼ
߆�OOs����	���n���M5�@�=?3Y�ӭ�&������kc 8<r��*�(:����Bvp��*�
7��혉�4����ަ!oX�is�Q�\�ا���n� t.��Ǟ.����z2�u�V{�Q���X�i����M��=�����,GD����d��PB�f��s'/��v�crjj��l�P{��������w�U����2��NF�1��Y)L_t?�69[ȕ;�`aDQ��:��G�^�����S��U�ݣ�*��P��dY��G>9��}�����>X/O�����͛����Tv� =�7�}o$]廃���W�B��w7��Y��> �|�n ��f�{
���v���������8aݞ������z=��0���b[�\�W}�1��b��L���_�߳k����QҐ��n����sb���X� Ot�^59����#]�T���߮�k'�|.[�uF���]u|����Ng�����Q�̕�},Ƥ��>&�������e�#�>�E�3*�^�-.|����/��6h�������OK�_���K�':�8���p�nڨ����Q�z�(�h)����!g�$+1ƷL�o�5�rot/ ��'[-�S���2Ja��y�<���XW�V���^�x��҇��q$�d� �=j4�|��-��|h=����c�����kjhl;d����CS��g"��D�_�/G�4=���j/�X0�(G^r��]5<l��~I�#�P�ipEiL�����'Q����/
2LM�����%_��C��OG�4����+��B����TM����P����_�p�a��!5�>�N�W�⿖��4@�.�󫈛j����Sm��?N�GQ._~�kyĲ�����p9Sd��N��?�U>]g��	E�(��dJ6$,��ǫ���/�m	#*Ar2����r%^����B���Ɍ>U�>)�Nr��� p�L�N�{��lrɖ*�����2 @
��d�F�qu����'{(���Y{ZW[�rL zr���b��t����:�D�"����t/л ,s`�6�#&�+=
φ��D�'ïuy){��0}��, ��WP��@��?wn9y�?�#8���/4� $M���{�/歎���eH����?�)��7x�޽�o���g�	O���z���+��S���䁐q
D݇wE�0x��NBp�!E�Y�O�c�N}:�E1�g�$��m�1͸5�
ޤ�Y���7.��Wl��&����W���D����������z�5	�c�m��1g�c}zi~>�~��t���ѕ/��{���Vo�D�K+����',z}�v?o��,bwdќ�N�Y=x4ǮI�le�4�5�~�����C��֏���11����;�s~����"��|n��J�� ed%�Sâ$/yO9n=y~ZF�X\I�齗k+�4-2!W$�´�A�V�G*~5�,cY��ݙ���{�*ġX�~�+�����G��3D\�P3�����/�$_'��#"8��q��� �i��ܰ� �1</@�VMc��~T��g��jy����'���g;Pa���Y��%�Z >30<��i5�����!kK���MUt�<�
�]������9�h��}
נW�8��qҖＫr�:�#5�Xb����pV�U?5i�ʔ,��e��c�y?�����}�ȉz�רZ�'�2ؒ��?S�
�BZ��w��q�߮�-U�(F�+aӶ�E��5&�����|��l~�M�Ǫ�vz�<ն���&��3>��
"��������D��p�a,v����iA|999p=_�/�B�,��- Ɏz����k����O\�ݧ��(����&�t�C5�A��%9fb\ae�d�������-�R���r���ѥ<:O�V�u��N�z"��}�	�*��bλQ:�.�����`ko����u> �s��u[�[�׏l��wg�MM�x��O{���YV���ވ��SfYw�P.�
�v�w�)њ-�ּ�z� �X9f"�:� Gc6��N�T��Z�-S��b_֠Aj;v��h�?�bH�B)D�`f�u�p���M���PT�D:DM1�7>(�z@��kX9�76�wjD?o������ԧkP�HxJZ�zݫ�%|w��g(S��O������x�}
4��#,|��@�`F��h�YW6"����Q:_�ji�!�ó54��l��;[�e5�j]<...��#S<<<�}�"9b�.f�]�#D�������1����(�O���OY������ƯS��7麸�u�6��#������S��)���F���Q�Ϟ��U����&�L;�̼u�/:^㼱y���jX7 ��,�X}�m�}����$�;��jm�X�s�8�����ln��'nSv^V@����vӧ��l��;Z�B+%���R��z���rX��C�����7��%���,��x�>Z�Y����A�bWۗ���2j]������k��rzw'�޸������x�\=�d˧F�3�s[t�tg�q���9n�,q����D��:�����M�l�_W�#�:��<��ӴD霹P��`2�u||iyYE�n�sI��Q2����H�+���:�nc{P��~RB0�w�<2=;?��?�U@'��s�m ��'ͦ���XQB �MTj�y���<;�s=��k���Ч��sP���v��%/���)�.ki��-��>��r��WZx��
Q0N�����=��J���zF��hԞ�|��ۭ����^@�6����O��a.��Ŭ��c1���{0;u�e�,���5����$���	��䋋�T;��n�]&-�*	�L�����ځ-�j\Ѫu�*�� @^��_�:��P�����I�xv�>Z���Ug2�l�f����/��Vu2�[8)�ql5����8XX��s?֤Bcj9կ�6s߆e��|�_��;������[�BH�Ȅ���!���e;�~��O&ޚ�;Y��c�����/?��퀯���{���Ѹ"����t@@�¿l�~ߙ�����i�P�ceXJ��$>K� �,~v�T������\�Nt5�m,�0��f���q"z,��X�K��J�y@���`��!�J����Aw���6��tt��,�j�Ƈ�ŋ�r�[i���zE�EnRw��P�D��=�����!_I�d"��T���""�<#��WBN��=Q�eN��X���YX̴7�}�@�*li��FQ�#��7Z�o���#��W�-�u,�S����D
�<�g�no��`�.�2�5���{R�T�V�~��9 �Pf��3B�L�}zz��qjq��p�>auJ�=����w8^�6�!�+8o���K��(Q��ag}R��hk���c�`Ϟ`�^�� ��Q>$0�*�>���:1AQ�W�q}}�x2�/>6��������8yT��୭���,<||��Ck2zUY�[��<U,F�q	�導��Ƴ��lܰ�.���RX��Y��<��`y*�RV���%��}"�D�׺�|��R�b���qcXl�-���k�w�bqryMMT@�;�,4�9QX��D��/��}��t�@m���˼O��s���&TP.oL)�a�C�;��h,�~�6�Fu
���&�.�/�O)�����؍��$�D_��cK�`���4S+0��y��Uf��Q���h�l���$�҅rĽ��uR�w���|B���lu�;�^.{@�p;�:E�?���i��V�ߌx�U�1������I��1�j�!�)�]�3���YP���#I�j��eNV��7�#�h��Ԏ�|���5��h�t����$�(a�u��Ky����`_SK�ʊMTL��r������p��r��lи,�_����F����YX|��87UU��Xk�gՌ����Ja�f��|���סMKy�������aT<�V�T�L�̞2ΏB�?���[���{�%�w��S`"*7��Y<��J� ��ayy����6y��/�)�ttt������:M�A/H}��G�T�����aU�x�*!C��X����
~-��pՄ�V�20d+�@O�Q\�M���C=�A��D�&�H(�&r Q�˽C�|��NH��7Yx�I�F�D��k�v��ז4���IDŭP}ʲ7x���`w7;��K��S��H"��|x#���N����$p[�o������b]�"N[Q?���Ґa�z����"���Taʜ!H.�[~�6Z��P�c�>5��m��E�Vu�5r�8����C���9o�����t�p���,���Z�>|�Lk���T+N������ؾ{SW � W�Sq��7�`[���6��r����N#n�ԱAඬ�`��.V��ÚĮ��>��g ڃ2~��f�U��lB�iM~�(<~`�#���<Ԡ��+A�C�
�2~�st���f,r�a�=gDi||m�f�;(Ң;F�f�=�~�K�9|5ۼ�Fb��Q�(������3K*�X��&���[�%˟g���U��#�-Ǜ���.w�R[�W�H座&��===��n����Z���Q���;t|��Xi�9��/�䲍�h���~���w���>%e�:8�ޤ��"a���S�
�u��5���WGK{gUXD��%��/�=z�M	i9Vҙ���P	ƻ�\A�搰n�k�>3k�rhXߤ���������;�V�*	F�����<���iI�䪢"�Uf�[OmV�1��k+%��Ye8��ȅ,������g�T�Uϝ��\�ŕ���f�:-(�s��(y�jN|������O�UΛ�b�4E�RE��em���0�VnK��ػ�s��=��S�ӛp'A���Qt�㭨��jِĘ�����;��_F�j,���C��{���;����N��^���^��
|�w��x���V0b��A=Ekձ%c�L�b��`�%318�����@m����i�B�%{�ZZ'ڠ�����̟��6o�����UNN�%s�J�[Z2��.-UӚǡx�P,�.�}��_��S��wA�pX6N䠡 ��$�V�;����q#f�%��n}C����.��ض��u���g���w��bi�jo3 �c����I��("�/@��s������6�^ŭ��8�"/eo�g6>Aa�7 ��ir ۃJ@� �d��_2J^_��]\h��v5���9}�	�{+D8y0��v��+k��YO�8@׾�ӾJ4	�u�&�I1~{����-��s ��y�U��C��\��@�T�J����3Ȏ����^��yE���L ��lP;�8���{�i��18��Ih��\�_y����DC��`c�7��<�����[��@G�򖊜2= vZ�N{�4���E#>�O�#�va	�ܜ��]�Ki�=+c�/����w���ވ��G�'�7[��
�{C���t�/��E\@>Ń&{yw/��j|�W�xL���ϴ�e���ǨY�P[;����Q�Lu8��A�C��/�Z�E��y.�,]��ea����Y�2n���Z��хU��/�Cn+���'��8e��m�A��3�F����IB����y�6�x3`� �;8SHw#���Y��Ǌ��� ��ʢ��<b$�At��2�K�!� ��D��OȥNt aNP?_~��qj;���d���Ťn�V�ex�A�Ņm��S�����j�s[��橚�� � ��n��=Vs�ws��Ǚ���$Z�K\^�[w����R�K5w����˼;a�vc�3zS�8�룺r�wZ]Q�A	�	���Os�L����U�q5�3i�h5��Ldx����G�ֺN.5���+�����ݠ  Z�Ƕ�ܷ@��SaS��ٸ���O_5��x�@�(s̻z������43�Z9J���+y�u�rBڻv>�/8�VDx�Iz僜�i0�r4��l_�c��0���WTV6�u}�H�R̪�wĿ���9<�����W����,�`$��'RI���1}p[h�UǙD�lg52U�JdMud98�t�	}�DQť�����ag�6Y'�+���P��d=��\��&����w�jp�=8��ź*?`���:v������t~go3=������=#��4>�mI-g��ӓ������>"·Ԇb�X>]��z�O[ ��!�M�f�"�����'��KX�I��u%U�'?=������V�t����d�
��ހ�a�~�����(���\`��l����IC
m./��ס��3>>��}�~����x�?5�.��S��8߉��8D�J�]�[��0"����/j�P�֟�돊����W���Z�TXi��Hs�w´�N�_����;u	�	��LLL�������
a�AT�/??�*���B��
�w������_D)2[��]Bf��>h3�ե�r�Ԣ�E����V���um�Qψ�vS��U]��i�KC�y&�5�� qͫ��" '�q{��@��o?+�Y	����8����#�'٦�ǲ�4�ػ����^/����.����3l|1��@�!�~����n޲�� R$�f���?c�}R��5�;�Yis�8e�݄M--� X�ˠ����6�>6��5�P�?r���S�<����d��p���N��H�U�Wc+[{b�2��߯�(M�^�Ri:��3KL��R^4�H͒���(�~�9B�aI(p�����wz�!w����4������ [!s��m�_$5M��Ѭ � }��QIĞ(|����g� ��|�p3yp��w������Ҭ�,#�E�dZo3A�ë'��e�֭�������lX姹d*�b�/�ܧ%ˁ=z�����;"I,b���*�����P�{�!��8��b���@���ǲ��w-��6%']�b�(#b�=�V���C0�����w�o6~kѭl��O���k����v��WVj����bU��Ѓ���q&� M�Ծq,,e���.�'��$+��6��CT\�¤�V��l�
m����Րq~[��6%�X~�I���d�/�hx�"�Z�t��{�y�2I����@Mw��J6A��'�����j��Z��p�)��)"��KF�[���;R$���X���ς��*U �&2���8�{��C�ZZ2RY��/߼���9=}lf2�)�r��tn���=G?�^�G������א�8K�2}�Zf��ld���X����"�2������S��wD��ˇ���T��k8�3�����cV�(����y{<p��s8Kj'E�p�e��G���7ԒW�TQ������<!b;���Ō�˩w8J���xv�g�Ծ}���?_L��;��Z��8I�;�bxz�ȥ���I	��	�(���k�)>^X
��6?������蜌jS�Z@��U��@3�!iN8$*��o��-+��\{�p�c�V���y��ț�6c�w�qO�^M��%���r� 1D�J��&3���^��i%<�:~,���"�.M�>�A䲬�|
�>~ȏh���7и3��jҼ�Q��|ںrm�!X�Tӹ�[qY���!�߽�� ��n!m�� ��ht>�'%�F�L������	�����:F������WxŪ*�N�+��D�e��VNn��WD?��M��ʪ��J,�W8v�=��ܓ�2��u��]��>`���6"F�&��l�=�xd�A3.���˚Q\$xd�
F��8x�__���}%L���H����Y�2�f�tq��J��GO(�/��L�$/'��ʞ��z{��v���z2=��wY0��)m�)�P�X����D
��.��?+�b$��~��������p���������K�ȭ��b��#�kh��[w3Z~��-i�-��V��{G&�4C�۱J���j{�*�NE��j_��2�t�V�XT����_���|n4��۞ڼ���Ӆ�w���@
T%e�@8��]��*(�Z��e�yYM��)`��I�r�8����Z��JX%�9���DGl�y짬��[������ʹ}���H-�m����ɷis��{܋�}�U%���}d@e�9��۱��XZ1��2�;���0�og�ķ2E"F��Ix}-�T����F���޳`3�B�֓WM�(�~������m�5}'����_�߱wO0qʓa5�	�nps��枞ׯ^�yq	{�X�|~	�U���J�h��V�f[���sa���w��y����]/���Oe���P3^(n�Ɍ��/�6�`�u����&X��g���)	���`�'�!����v��IMg�$����	�5����O-l�R��U��1��f>�Q�w������V��f���`)���`�&�����v�#�q
����Y1��,z}W�I�.�m�Ky���?l���*2 V�֣Lx#s���@��~5�v�W)DFG�GH��H�_y��L��ޟ�kq�=��p��[[Г��>Z	>�;<`��d��"e��|V,�y�B!Xې!�Q���>l�}ơ����,�l�uܟW��2��� �"��E&ZSb�/�o��V�9}%�Q���S�����Lq�����t�@��1/L�:D,� eߵ��|���YZ��f���|�_��9�����;7���zn�~5jN�0_'�b
5K����i����T{�0b�o��v��@�*TB�,�1��2:��=��hɯ_�x��5��(I��zg	�?�ZS��l�4�j��Z�ɗ��[����d�1�8)f���7��?�R�r>��=ف��3)���������\��W��`���Ad������w��/��w]�/:���għݼu�B{��w6c��Hr���>�*����}��$s�ٗ"��{ϣ�4��@��lFF(�k�Y�D��u�s�\v��fZBl�Sm�wpA=Ϸ���l�g�hOо!��Q������)�����I���*H�������D�i��]�!�хO心��F��p
i�� a�D�W,B����P����2��Q���R��Q�~d~{�e�R�Я�'�ML1���-��z����؝4E�D���(T@J�<v��<f��#��{�kr�mK�e���&��%�4�w�%�"���	�F��M"r�T�gxʸ�?|ѣ�3���Z9���a��.�b�U\��������~J.� 9*g�y��q6��K����U��2��&�G���9biho�����?%���!^Aˇ����^����lu�4�YO`�����O��
x��������ۮ�:󛗟�2�ajR9�ͳ���%�
��SL�������Ir��k"Yc��\���`6~����κ�U	�,4�ʆ�c���s����d_���M��|�����X��/�J���բD�y�7���۸ﴩ���أ�Lux��������x�2��l�j{^������(<��R�@M{�a�QR�/z����l~�|�6�����>D�	Nb@JO��r�ui����S��Ə�P������<�&��oL0���I0}���>{�U���K��31�_@�3ʓ�v��-I�%�#6+���&�U��j���a��/��\�*���J����m��\t��T&��㏱pL�vrc;�Y;���#�c�2Sm���o ض�K�����a���"v`=�=p�7���� 8+~~�z=��V�А�a63P�yM�sq(��ny�Z�����=;i��[�?�����Q���h3����q���Y���y��$l�֔��_��L�.�D��M� 15�ڽ���bd�ǿI(�^�#�����\u�e]9xr�0j�3��LG�Qb^�
ݤ�dt�ʞ=(������&O@�==�߳�`e��?u�mߛ��~�iCL�}A݆!��҂�Q��	*$êߵ_LX��4��6r���Ծj�����H��o
�խ��6! �*#� �N�5%WM ��	�
���_w�/ہ���f.'G��|ZBhj���������P��x����{�ygۤY��{�G��he��Pr�^�	AKK�q/�*x��I��^++㶟f���H�;�Z��f笭���_���Q6�����3D�'�8�KR��X�4ʛy�CNi�wEE	�(�x��>ʅW�����t� ]q�]�JR�ۺ�"��qk���-���f�<�dg�j���?����4˗�R�n�?UA}{W�p����(��o�����?��F|+`DRs~�o�X���;=��k��+�?M|a�DGVf$^�\�`�=��0,�%l wQ��b���Qr��-[h,�!�����������-I9@~�­<'��\��xț��ar������"��G`[�W~)GzFF�� �/��qO�^L���_bk��&�
�������H�Fx_��]�i��9	��}ۯ9�c�c�pK��@={�8��K����~��v��qƼ�ֺ�Ož���-|Q�a��~qʭ�6������df~�A��^��mR�rQOՙs���'��x�<�!�f��ID��<]ӯ����tB��nq��Ч88��i���S��$ �2SR(Q�6s�p��u� ���Đ���S����yp;hI��ܩ!��X�U\p�ξb��og����c��l����1�J�8���W�Y�@�Λ������/ځ�Y�b���VdBz��h�,�HX
�B�/����QY��+�=��t�K��tUܟ��&^i�ݣ�j�.{�T��b7�	�}����O���N-,v�z^��u���u6���:z�ôs�����A&�ǆw�%�YIqV��=.0���(�� g��|�����a��foCO
=X2C�5ɚ�2�YP����(�Vh�/��$���!�!G+�1@(C���9oX�n��:ID)Iæ���X�D=�m|\�����s0�2|Z�� w���J�p�a����� �(:..._�k���̓�j�]e���W��Nt�t�p�P��?�����Bi�S^�0�Fr�d�y<p���a���Zn�X�*,J�����ʕ�T��?�O���y��1��+Iw�j�ņ���?��>�եd����WUou|�ۓ?��p����)�!�l��1N��o�\��)1�m�M=�±���ò�4�����Gp�\�@a
�i-��|���PxӨ�c˴x�O���-�-�7�^=5%~.���	/�QW�M}���	i	�����ZD�缆
-e%�C�m2C�ƺ���6]
�<_�J��ň��oU��@�b ����ye�G#/����mP���E:bø��L��S�x�1�e��is2A�s�U���C�@	j�vɺ�xu ��1T�E�E�5�����$����$(5A�؅����������������p5M����,ȏ۪^8��h:q�:Y��&� ����b*�{��Sw��xCju�xC� 8�N�=����SO��������1p�S���,��G��6~J��V�k>m���&9���ZTbF�2�2�V%miQ䖼����Z	}�x4i-�����I���8W�3�&���U��z$Qh�7�����TY��n�Q�"��<��Yl�A��G��M�l��_m
o~� ��&������<�4�����	U[]�G�_$g|E\���EܚF����*6c#%�)o~��f��a���l�7Aԋ҆������r������̗�@�=�Ç>qj�+I���M1YK���W#ÉG��
��m�&k,�9n�9����5��v��X��"R^hԷ�v|y)���:�>+�R����A��=��������y���z���J�y.�����0Q~$�s�����>L�F/`�!���l�E2���ѺJ�JEӌ�Cǩe�����D��$8:�����͘]Kz0~�)��Ŭ��?�����u=��CW2�ه��G7���Gϰ6�/�o>��]��j��%��j5��F�M����]�.��$�u֠��c�����K����j�7�2#'٢���LIK?��g���.��@�ՒZ���c�5�G�HV�J't��ilF4i��� �5�����S^B'�D��/Bìv����'� ,���m&��m�C7�9mgy�X �S�Qh�p|���v���쬫G-���X5Ҝ�5G���$��2���D�l����}���)$�Ȳ�Y�\;�(�p:��(�I�zx�;d���<N>ȋ�j\}�_<}�z����kQl�8e{eu���!��5�$�׻E�9A�D�����j�^λ$��O-�t�܅<x��˜y�~���R��[\c#��abܧ���+42���J��/$��f��<P4�e���\�8ON?j��S�3*����5׳���z�˲�kNpCQCC�Wlu�@�/Er�U�p�l�lAf��SEd�o��f�q}<����H&ِ�Y�6��~i����mg����	-:_w})I���dH1i|].>'��h�L~<�x�J��� ��UBv�.���z�1J��q��]t4N��q����v��'�q�ol<�Ȕ�@�v����^s�<Ӫ�KM��-��2@t���[8/n���H`鄑8j%�З����(��]��P̖d��ِ$1��U3[M�"���<�R�"Dr��}��I�u��]:���\1��%���1���sP�Z���� -ʘ�Hw_̼�tZ��|�Wj57� ������ ��M5%�BP��s�M+��&΀�)����V�S���=��a�R�{`i)�ŝ��-:^O'�u��?�[WGfhh�4(�ؘ�4�ǣ1��{�e��W�Ѵ�&c�Ke�i�D��'���Wa?��_�(`9IczȾ�V��1)�L\�B!���*snQ��>h��a�]cJRkE�Pي�D?�˦�ٙ�VQ��>=L��7�W[���9���!6Wz���'�Z�wM(�j�7s�MٕRY0��6|:9p�Y|��O%?n���Jg���i>��<���zB/Y��J%�,�缁;r�9�y%[=;��~���῍:��5���I�|����A@��p�����AnP�<�R5(���͓�G��.\S�y�H�f@�����L9I��8;94�$��ˁ�Vz|y��r������v�	��=�L?�cυ� �Fi˨���^x34j^@�o��!�G�j�	E��Ȣ,��*VV�N��z���q9'�(DL*��v'X�CJ�T��G��SW���Ō���U���+6Y����[7K��>���k�iT� S��t{9\�����^�r��r�0"Q�!����ͧ�$l.��3�E��k���	/t�2��"���a���d�`z����mL��(�{gW��~�l$����>Zխs�U,���(�5MQ��g��wy�q�E)������F��Mt��U��|����I\پE
�	L����N�zB�{��n������C�c�M.;����/S;;<p��1)|6<��%:py48F961�FL�~]8j3��փqW˪`�|NTggKv�T�2^=�8=����������Z���i%$�c���G��v=�zihq	;�k� hs��ݚWE�S��5����\?>v�q�҆�����J�*��(�"��������C��3u���|���!�/)�5�q	��[��VJwf�s1�1�,��d~��Y
پI`��2�_M�Z7���!7m��V;��%�F�m/�G�0{����L[��@���{��;ѕ�3��̵+7����vA'8��'ײ��>����4�� }V�RC"gjH%~��[c!�nX�xρ���q��B�3�n����̺�ϐ
��;�n�i�1�E\�����I�ͧ֑��@l��^��	����L�I��88�[V��l�r�]�BZ�.�*C�h��gK�6Yn��,:���O��=���l��\<F5�)�=�g� s�����3:8}6O=���N��?&՗�����*,Ϳ�lӪ&��I�Ƽ!��|ꑒ�W���I�*J94OS���.d�R�5m��{Lo�;�h��X�,#)M*i�i��F�頛A�F������Xl},ON��l⭁��Ėo�z�a,0�1��/m\�����<]��6i���.���}��d��.F�&팸:�\���*	J<�-��7��D}�R���$)�A6�FM���u%����Ew��.��+��eO�:�&�V�OjQ���=O~���9n�Y1A�x�R��/2�l���ُJ�Fڝ���$Ɲ�;��;�g���A!���q.
E=�A\Ҕ��(�mp������٘�m嚻���4�_ȥf�/F�jx+�����\�졿�nа�����6���C�#�<���v�ZX��ɯ���U���l����D#�g����i`I[f^ףl�=%�Ɍ2a�_k%�ӫc��ݬ�mY܅'=����߼T)ר�0���9�yg�����%/9����%d��*���7�no��/jrVA}4������V�e;lHu�����1L%z���$��E%ߝ,5�bU��[�T ����c�~%���-c�c=Q"��8):��ğ?u3��AA�f���⦿Y��9��Z�Nt��5�|��8/��
CJJJ�'�7$Ǯ��E?��ywV0�e1I;+�I	��V�^����{�5<���Qy���a�=�Fd/��o��Vv���|�1��xo𔺯P��Q���L����y+D]^��-��^��S���V��k�:̅��ւ���l�`{k�h"�T��@> @�UP�XW����G{:���#�3WG�Y���{p8O��K��?�+�W�R5̻��;�X��-�X��_���Z�i*���ݝ����jqn%���	('.��M��2���FC��FÐ�u.���rt9��ye"W�:p�
�UP��~w��Ck����VB
_Ϧ߅�
?�B�m�eQ�0R4���r�,_���@2��S����}G5\לM�1>F����6����X��6ʁ��V�w'�M���z_�n���i7������n���Sb�����n�Ut�jX��1F;���b�����|��n��]�s���&�)U��piƬ�����YB����k~�����<υ"�L�����ԇc:�}#-�d6ߴ����fv�h���ܹ�Ff�P�HǑy�v=��S���h[��3uR*-�����i�J��5r�J�}D'�	���d/u/�j����(��v���3dد�ã��˓�[�*u'^���2,���A@J����	����$��n��e���A������������.x�㬵�>k��z~��yI	��C�iD�RY$�bu��ܜ/"�/����Z��e�o�қ�lM>l^i�,�ޫI>�ն�+�ǭ�����������6�j��o<=?����\���dp^��쑖Ο��]]�0���T�z"D���|pP�����5�^��{w㔜�6�@��8_T��
�����=<��p�f/����u��;�U�Cv�l��\3:cxؘ&�B�;��͑��������na9ws�qG���J��bٛ�e��n�0/�(�dqG��H�`iǐK�n�����p��Y�I�L�XV�2�}�0x�Nm<�.rx�O;G��;�j�!"!�k+�~݂�0��xU"Y�E3�kx��81���ȃɹ,"
m톶B�1���C��s]�j�|,dh([��<�:�7QV�CQ�k��+g�$O'�.*jy�]�1�t�1	�_x��߇p��y5�[�Հ{G��z���|7�oC���!�4����C�H,�a�kļ�V��3[*��J��~��3a&�����7s3��
w���җf[�!��YL��kD����ܛW����i)�!0�r��is\pMNE���gjP�ýV�7�}�U�|�]��j��&�m�˰`��u�X�ڱ�G>Rz+�Fc'8ϊ�:s+ۛ<�8p�9A��ڛ(���Af��畾CeY�zw� 0F^�4|�N�{�y�T*qlr�%{�V�q)�:�(=����yzg�F�G��kJ�P��K�>�v�4Xd��e`}6X�Ou�7��g���7�VĄ�����&=�7�����K����<!�'5�a��¤���o ,]�����C���3s#���7�{i*���� b���[b���o���hW��PZ��_G\#&�̺��_�/���mh�6�k�}�	�7g���`x!Т2�Hj��!��൤��m��+^O ��E��$�y@@@���F��y�ݟ�rQ>�hiko��Nԉ"��<�����R������0[�;0t:�����ygR�,��W)J�rka�?�lq���+��������T��"9����o���xB��j�sG����ׇWs��U�4���HJ&��E���:�E����w3�#�c�YK-d9j1�S|��[g�J�w�֏�t��!S&�.H{5�'(�"�r=��D���!��4po���͇�=�]�q��13�aA\��.�;�����>�'�e�k뙧�� ��uE['���7
B�X�"Ja�3�1b�pfWB�p��p����Aw��rS�k"�˽�$��r��;^�Bu�2��h��f�D��ui��~��C�B�YI�i��@
# /Evx��Z߰WlӪ��=X&|���d |4���9�$U���W�Zi�����I��y|� ����pv��,�0h8�n�.��n<d)ȿ�����yJ@J�)Db��lw����o{˪tX�8\|��C������4A\c�����Dm%H�Û��%�y�*�<ǌ�<*`�K&�~��y���L���Q���j�����|*iG�<��H��E"%8�����C���	�	��G[y�V��C�����,P����4�O#~C^�(�7��h�q���Z���a�I�)�(������c����ɼ�ɨ��-�W��pW����ڊ�_g��2r���|�� �*[�����7f�c��Y2��e����If�c���T�-�;
ƛf{2���/��2�-���yuY<,�Y՘�1B�3,��y+`�	�e������;/�xx�N3ws���h��B�,i��c�\�;;�&! ᇱ{�GS����[�j|u�Gǚk�};�ܦ�<O�
�F���=vRh�)��M��ᱚX�kҟc��PжR�CKn�2θ/�Q@#}n��23�[�G���A��68��b��L_����Ӫ��d-5�A�2�	�Tϵ߿��ՖK>V~LđQJ����<9�*{�^��|_]UQQ�%�� �0���Y��'{)������Op:�����<�����ú��y±��)�W;��Î_#Tn�:Z��t�
Uh�I��"+������j��$LZ���\j��� ����	��?Ə�9�kMn_�P�+k�^<�r,M�]�_@PoB��qR�DA�b<�`*Lb&|?00�<H�^?H����k���h�:\9�k�e�����z����p���M�Q�����v�ͥ����Oz�K�ٺ��m�׆o� c�$�AdS'��qӰ�&��X:,�o�A�IfM�F�-������%�,�S�!�`����0T�T�Y��D(���'�!��S��ي�)y+�gA��ݖ����hH!�ċ����Ra��h����$P�?C~���Z	DX)w" %��N�*��H<3n�A��11nƑ��k9��[P0��$Μ����#I�]vHcӳ��a�����X���E���<����9 K�U��I���r!ޔH��n�4�+S@��7^?�q� �6L����3��p��ǌ�q��aG���F=a�r߲��2]ei�ql�1s�	����v�>��"���s#� � �,�YYs���������dU"�Wo[���WRq�L%$n�6��xt2��$%#no�`N�yq�!<�Z&z�6A,���jc���
�%��+crAf��V'�͢^j<�e=��_���P�Ǵ�B:���d���?��o"1�/q��q��ҹb��kJ���{$V��ͫ(z����'O�J�M�[��*'4Ī�� ��� Q�BlT�i�5���Ս4C���+��a�>�k�"���S�P��ZւQ�j���Q��y{"�����w	�B���n������SOS�(SJXE?��iy3r3���3�a8���?NQ(�ԝ(�YW���������"x㹡�Y��G;[�F�y�~$Q�4�5[<��^����'�������ٽ��S���x�S�����K}���X�����܁�N�;\��:��a�#����<-M��,�E�^���^��Z0T�����= ��ZZ�����֘rYE�cȨ����&������@4����������;� �p]���oL�6�8�q4�414"��\y�<6k��yjzm���Jy�~6��C[��B��~�8����ʸ���{�:o$�1~��k���®�D2�����!jV)��Z;�KNX��Vȼ��x+��V�)���� ���,� >���뵄�����(!�� |��u���%��?����^��¸�6��P �ڋ)4Ԭ������)zªG>JL�SR{\{V�2+�~,)9�65��{��W �lEUU��"Τ�椮wt���H���Ep�cZ����z���f�o�+�O�9�\+�ΎEI}�>O�'�e*�ij��Q�P��Km�� KZf'5�ہ�'���π�/z]-�4R`	m��뛟e�b>�'��a��|$�u{�X/m��,A>�z>���f�<ޟ|���{;tN� 	����Jf�ۤ��UV�,�窫���<� �NkV��I �5�E��,Ņ����x*YR�2`vG�����me��k���0��~ٛ����-�S�f7K:5o��[�:��>8���p#K��\���~k�L��\w�1��
�����4��$�|q��D�S��2���m�o�TaNE%k��]�eҀc+�o/*�]#sSѣ��tF�WO��<�&��b�>�av}���<��R��E�T����q4b�;<P�ԉY���97K]p�e�o�_s-T�c	�}��%��b��8����,j����z\�?<�?�����y ���sv�"�b���;�8���;5Z���a�w*�f0���"#/��8
�A�'�
	�{���4
�������-:��I���d�(��M�]�ɦ]h�Q��-S8~u�(���ʓ��Y[����Z�L�"o���I��w���ʾ.`ބ_c�>Q���L6��!�c�B��+��3Ǳe�d��w�4��Z�Z?'�3[�Ωab�j�zQ˄��d����>�gK�43ߥ�~n����d��OLrk�(��ȫ��I��ׇ�?�"������y��x	�;��۵tXt���f���$<�D$|��s(�f����v�roez���)z���Sv^�败�ʗpv��=���+�%��ǭ�h�KLu��c������� Gw���YB��|*
��N�ҍ������q˻�S�M��n�dٜ;0�P���;�:o��9��<��*�Zy�:<��?�1����H�Y����mM'w�����2R�D{�u#����\������B��n�w)�zY�/bu�3_�Uy79'�{ﶪ���Rc���������[Φ8rb�$���'W�~����P��q.*R�����c�ڳ�G����Z��2h#Y�����=��T+�Õ(=a��kzrA#	\�@!�z�[|�^�60��~��a�f�"hL��R��o�����>VTT(f�	�J�m�B��yr�/�\w���i���G c��nC׈���ν�M���B{��X��ޯM}j\2S����ٿ��_�kcd�:��g��ml���S����T���qS*G�v*Q�j���]�q��uY�;u A? �O6kDA�j��ﾉ�d���q�A7�<�ڜ�Ja�����V�i�Y�Z�:�]��+�S:��Ӊ5U��S�B��q[l�Ta~���B�S��_�n����|��5cK����j ���f/  �5���3ı��;W��ؘF攽��_������YX�d��"�˸.g^��n����ŋ�{����{F����xi|�Ъ��m79ظbXo��V#W�����1^�=x�ΰ�N���O?uu�C �2&-��1�i�c�c��Ăoo7����!UUU�Qr~-�_)9����s|�"zᣅ�
f~g1&r\D��_��ߥ�w���GC�'02�iǽ�^��K�ra��Ҏ7+q"W}�m*�@D_DF`_�S �si�J��R%���Ɖ}�,��e��u�n^�G/�åN��d7Oם	r4�tq�}�j�M��­�0��-�I�����7lQ5�u���D��lGD��2�p_�0r�Kԯ�+��f�Q�e9�v�-œ	m�6��B�����/��q����ty�\d�Qo���D�r���s�$��ڔ��@���6	~������Oh�Wh4�(��0С��}'31L�깋�����[3�,ֽ׷�O��Sb��
�m-��B���O�||����g�2tL0b&j������f:ݲ�۲�o������o�"G?
ƅ_T� �_^!�P�h���S���>������ήO�Ϩܡ!.\�2|�+��(�����46�k�⦻���l�vG�VF��0ț��gu1�^��0%BR��W<ؿ6�ݢ!��OM��L���J�)΀�.V���������A�'�� 9� ʇu��!��\Z�Z�'N�.�$p�遧��Mmq��}��U��"��i�֜_2�6�ܓ�x�,���C��?���U���������V��Y�2�K<��NM ?���.\g���7��R�Q��v��h��呭���Z$ֿ����un��[W���@��T�q�|���-��=k)�C*�|���")�G��Y���9�3n��z�$x���D�o�\�]e��fQ\L�g.�}���(�������k6A��R�ǝ� ��ϭ�$���hVu�&��V�#�	��A=yh��`�C�/а�����o&��-�!��b2�Ȱd�x�.!hJ���o�ı~���nL�hg����sQ���O�k)�j���>\�b�lki
+K�٫~L/��2T���=��Ǘ2����ug�Х��6-q�� go^��A��@/����q�9�2_���f�Ӳ�� �ji��u��v3�=���J���Np�����-c6�K3�_t����R��-�c�����7FU���Eh��K:��G4זS,F����DE:�a�3a�#74��}�b&qR�N82�š ����?D�wR�&g��-;;C���p�e�h�2vgg�V�"l�>Ss���s�S�r�y�K� ��:B�����R�ps�Z������!��_ݽQmQ*����u�����Qoc�J�e"�(k�d%���r�����Z[[3x�������r4쮞��D��S���I<[�e�d�1���������SD1l�LΌ}�
�|c�d��˗��Zz����	?�r�<׸�/o^��c�r�F���f@`�Bg�$*�[>#e{�,��"��U��Q�#�5��"�5Z@˓ �`�k㘽%�NБą�cS��N��[��4��|����>X\{7�D;%��8W4?������/���B@�psC�A}��7�������"�N����_I"x�yP�>��!1�������ڻ}JN�؟�ڐo:S#�u<�ӈ�h�ϵvv;�L}�Bծ�66B���k�4P$~�E+zM����9�2�f���pX�CW���V���q�����gX�����NEnw����90^��1�2P-�x����Q�8H��ژ):������bǉ��;sw�^"a��ʨ�Xm���-ʳ~� �GB���.���d/�)|��I��w�}h�gr�g�KF��;��=��t�v��ţ4�W����DI�B��,jN��B��Y��Lmv���kd�=�W��T<C"���/���@�# -�y8���1su���t7R�8�+�����{W������,�,��H'�:ﷻ��w.\��m%�a�T����g��n��1{�f�{I��v�7�^���}^�z|*& �t$����hko�;����bἎ�����Z^�c�,������f�'��� �*�7,�d��)�!��$�@b�j�hp��L{�#Xkldw3���$�..^W�C��L��e�S4�h���	�����{�>4�gS|�SN�M�{W�ۯ�[z,�[��8M�a���>���2�si��F��.v���T�5����$V�k��a�G�=[���͍��B���V����V!G�W�؛��e�a|�!�X6!l�����}�"���!�hgWU�M��L�-:��F���>�0���t�2��~ReEA��|��C�w������:��!+�qރ]6Q���Jn-:�2:�1��xa����5xm�R�R���_�/ϕ����St��W.��G���֭r�_�quD��u���`)/�A�����ۘa)�I���������i<��q���
��e>i��rvs]�P񥺷L���(�:����3��B.�������T��ܒ�	������0�����`�~�˼�S4dG�5�!��f�b�{��ƈi�r�?B�ܳ��6_����4�{r��;,.r�sw�I�K=OѦCb��E$(�&�GT�Æ+n!�dF%'�ߋ6�L�<���gӬ�ޟPUR����򰯷^�G��I��1�<���a�X��>$g����rww�o'����SV��½nlM�~I��_�5*&��9m'�{��C��|~#I4V�'P|�J�G�'Bū*�&'��͞�ݱ�,����%��G--�Uv��PL�~B���a%�&�� �,A �h�EԷ���h_g�MKT�ط�:������`)����Q��l�b�k��HdT�+1@|��~��"��c�}(�S5�����ڷ��>�n�\�7�� �HI�G��{���ú�SJ�'u���gJ�.а�����VZs�Ke�)�/�S�x�_�s�ׯ�~��c�pcL�ٺ�\�:���!��%�ʋQ�@ޯ(+�����V�<�����V���f#����귡Ǹ�l�nlX�l��lᴗ�Ƿ��BB�����{"X_��X�T/'����Q��DW) �O@��H�4�^�0`�h 
�^Gou�P�6�߾�@�9f�[ў��(Híp�&���xt2�b�>Nrņ�`�������m�k+"`h:�g��{����)^��w���w:
^B��?�0�M��K��0M���r����z#�)���ڢ
�z����c7@*a(�� ��K�A!Jȴ��x�W��w��M�}�ABѻKP�C�r�������*�{���5Ӂ�J������ی���"V��;?6^^.�$��;vgz��X�/I ƣ� ����Ԑ�f��q7|�|jRy.P��}[�{/r���(�p�];�ܓ6$�	q"gK3,<T�0����7�;0m�u��_�
�ȇ/",����N�l0�0:k����;q\Ee;��1cotɩ�L'���[��.I�8o��j�݀���#��� �h��i��@-���y�>K�}g�D}��Yʟ>\LZ��"��/�;T��ϊ.ERC��&r�M�-Z����O\���uAc�c��:�U�fNО �jɔ�W�P�~7��������++� {��gS�ѥ��s'S�hX7q�s�ѷc6D߲��(�뭇��A�Q`*�Ok^����.�����!O��2b����<�)��U��X��#����|��|��e�@k�C���ڏW�C��X�/���ΎM����`f'BB{{�Gg��]at��qk�.؉}��~pX��q�s��B�] M&��Zo��;B�[0�Z�\;�nDo�#���E4��T�Z!� zS5� (W����ݽ1�{s�
p������_���yQ���;�1Ҫ�fqM��3|��+y��c�fs������NMc&;On��_	B>��sc7�T�VJ/�5����zD��f[yw/I�����9dd}S]/1^�t��8������g��6?�1���8�b�?�2�Fp�l�V�$*JI?��SW>�@ݶ1^��~O���q~c�Px ��ʲR&HT�GN����vbS�8~�^��qBH�qr3Il�B(��"���޲��u�w#���mO�E�P��� �å)P ����׃�?VgR/�j����d��`�/����Fr.cC�3�d�V��~��}���/�8��=P��g�qQ��k`f���<�Fw�1@.������m���  �<��'y;#��k��.�L�����U̵�UضC�t�v�_/�j�XTG+�c���^4���ͮ8-��o�� ��ST�y7(i��̇r!�R ;A@�E$���w��W[)��^����9�f��Þc�,,~�߬G)�>h�yO����A���-+��D	ģC9�l�9��!���/�V�I�vq⦩��$ߥ_�ŕ�fT�-�R֔iJJ���M-lP�@�AF�M/IU�[/����ҡ����M4x�\U�x:_�&c��6�+	���VX-��<�厅A�����ֳm|&L}4h���0����ȿ�7@����.�~�0z��ɸ�-��}�#��S�k!D���U�A�G�^��$D{_���W���<Xm�=d_����YsYQHdx����v�&�<���1mX3�=r�'ԍ�������@��@�=,O�����`��l��&[��7��\�����+�����M��X��k������W#���ND�{��O��P����7&DO���p9�������M�"���$Cy�o�m�Rubw*�f����O�Rn����z�nY�-���&w9�A�3�r��_�<�gf��Ty�"�=n!�N�Q=��d�:2�����5[��9I���Z�&����h� į6�s�M�:`!v��� ��{Yr|v�#'�pq}�E
7��3�z��tE���^x	�L2�~�,���k��Z3Q�(�����->�,[�0���,��Ib�׭jq��yvb�,��
�rkX�r�x#���z���e�jKɉ��l>)Qd$��~�]�rp�	dd}�s4d#�Oe��`)A�@'��t��B%K��d��������,N���e����%��ϴ�O3(�~��Bm��ײ[������ʏ���5Y�x�J��=�9<��sk�h�9�)Sx5�7{�C�9�]�ő 'NS��O.�g�/Ц~F��i�2��%���Upv^C� ;���a�k�
��6C[����}���od^|=��m)_-G�[���ԍ��Y��� �7~Y�vNտ�mՀ��X���cW����
�L���Y����FR1���b��b�q+C�?k>�$q�������4��si�E'��g�t�q�:*��8/��vYEMU_ki]a19��6�JW�b0:���b��w�S����;�!٪�9�ا�$C��Y��1P��L
�� �fd�VI��7^!�t`pc���!�jf*������WjOS�7��|7���ķu��2�� }����qMg% 9���4BZ�
������+~SD������k51D�4��W���&Uo�Z�K�;U��4�^_�C��=%I�]���9��5�OO �N�X�A����y�y�[�=�B��E�'�|5���J����O�u
uN��l]\��Y�p�܆�~)�W���C����;g�?�d����Ӥ��o�1�����qۏM��ͣ!�mϵ?ݢ�c�e���յ
HT"��*�B���Q���FJ-�ӵ1�N��#��� fc�?�(�9��ΐ��2Z� �,αςxˍ���2̽E�|�0 ��D��`�1j�Z�y���Į���=O`�seU��ҫ�:`�O�^SZP� ��Ce~�W쵹��`���M�����M���\o	^�'u��#M��p��ó�%�?��W���3^�SL��~���Ϋza$�d��zv�ʪ�X��^g�*/��$� kv�#s��"{����Jѻ���I�Wº1�3�d����x�U�w��*.|��Bճ�����	��e�7"��G��q��wK��b^�y�g�1^9r3r�?����QϿ7���N���R��Ԕh(2w�\+�Μ�l>�OI��a�wY�?U�;�R4ZΝw����ү�;����^w~��j����ZS!5�;�k���Ǣ���&.�6�P6�+�
|���:ZY�w��&��zج����MT�mrn��Y����?7M����E�M�/��~K"~X��8�"mx������k*g��~�~+�����^*m�#��,�pc3x�抓?��\��(KC:2L�\�"ٗ�&	�x��_��'�5�͈�_�ըB�㊘l�W�wg�BܰI(����Z���t�;��I��~�W.�Jb r`���JQ��H��^#�����A�ǻ����%\�'ܾ�,��b�6U.��uD�ǝ�g,!�G:ӓ�/���.��se/11Zǃ�1Tw�F~uPy:��H��9�;m�{#�����w��cc���(�je9�����Ɋ(�~{bh��1�3,1�(�N��d�JV�#伎;��i��@�
��M��c�`9���8�ٌ�*�.m�}���I��*��P�~��q2gex����l���������C�\�!��x� Xp�� E�Sp����q�����Z9���&�hW�_7�.&.���`揁��&�/%,^|��"���Ûw8��!�Dԭ�Ж��Ϣ �f��:��w��/�Y�
0��>�%���@�F�W��|w0Sto��bd����U�Qb�������N���F{B�����4D�6�"�੶�ٓ�"�W�Z�m���b�޸�v挿��w�����E9@�n��9�͔�A[8
r��&��fdl��I�Z��Z�5�Z��jj��*{�ε��am�^��H<*�Ύ[-NT�F}]U#;���2� C����(�]�z�@�W�[��MPT$�9��1��
s��1�i����?���w�� �J^��Օ��9��۔�:����%�2���C��F�d~=����QF�FE'- ҉�2��&nw3(�����P,Ρ'��Z�v��%���/�F:!3�B���]^���l� -�002H)
�Fs�IՁ7�6���AA��ͥt�M&�z��g�L¶$�����σ��Y�m�I��%?�t�ߕ�זFG���'����Z1s�
Q׈s��Ÿz�n��+"�W�E*�uSN�1���S�>���X���gѬ2���_��=Y��τe"�W�����G�p�Y��]�����I)Nr�:S�(g'�7����I��v����)���y��E����nN�pZ��?�D)���kخ��p4:���TZ�'!�3)^s
���z�(��H�$;������4ڊ;mȁaͥDR3��a�\����yU�=4�	�_�;��I���EUb�����ԏ������#��p3�0ȹ��0��������O#-֠��`	V_Ԅ@Ehv =6�:�f��p�9W�ܑә���o�s���G"��ɨ[�_V�^�3���q�^ܜ���ZZ�RWzzB:o=���o��3��=��s�6r&[��	_J���vu%�_�!���x)3��,����Ah��J܊�L�)-��+�p���'�}i�:� ~��0Qd0u��<SK�_�Z��SA�[.������[�"y/K�����̷ii#�vӐ�e"V��U�!j�b�)���2]��~��=K�tE�����U_Nܗ����o ��_L"�jUkV�)����P�D1����=�_�	��$��Rm���<X[[���ʔ��9��'\�z���S����z|+CU�S�o~iS3��ia�O�p��V^��B��x]�(����)��ʏP���z�q��[���+�}D5#�v������Y�T;�K0��-'�2�l+��̻!P%)�oDP�{B��҂i���ɗ�"?Z*I����ň�u����E��:�-�@��C	�H�:�,���D�1��s%�y�l0�|��o��<�%����9w�y�B��I{z����J�o�[�<hg���"|Cq��Zr�f��~ZQ��� $�nĮ�� �m�������[$�MEQ�^��6?�}�o�I�aW�۰<T�`Q�ݭ����M�L��p�2����ͬ�	-ނ[7UQ�v�-��\nߔ;�5�W��a��`a�8�PL0���y���ֳb�5"3���(=崋uc��`qL�*�	Οͺl�p�Q�6*�́�lqq9)��JE�y���ZX�0
 =�xB�:$�ĝ�xyy8㰙/..�/&D��Ue��nS�{��O�Ue�/m
ѾW��ͳv0\�\d��?�4A&�^�k�9l���g��I�y�3φ�����CT,,,%�U�ԕ�n�>JV0�ݳ�n���e:�Eʽ�=���0X�_�f}��g�yߖ{9ݎ<v�]<�����Ł6�0ʌ��7v�W��Ύ
�㙆�+���F�@ddwǦ������tj����%�!ؗ����e�,�ɓ�W+�{��lx���ht/��J��~8�	�_�ۜ��60���{�2?n>q�7�w�wR>��D���?}�|D`�?o:�=����{A���9�t�յ�h����"�;9�%D4ז����Yu�?S|\2Y�Ũ]��y�ͻ�*1ۂ&)9������[��h��]��|9hf߱v�Mf�8�[����l�Լ2G��S�P���NEe�j���׀KVl�x�`i�#O�@ET�;-���L�f��֛2���3����l�B���v�m�_�	����y�'��o��}��P���&�Awy����qj~���M��������m�{�����׳G|{.|+Z��j�4��ןx��>\�Fx��A,:�#���>e��v"��n�FvW�ju)*��K��& ���`��S�k���zy���$Ņ��ԕ���ӱ��k��=!�h--~2x2�Z5'h����V�kgGO�|�M �t���X�d�,��Tu�����9+N�����c���,�����h��g�2�i�`	sc-�N}���\��=xk-bo��BY����*�M۵�j�uN �]y���o�В��L�����-�i�]U�/�`.�}K��gR�\�Yk���7_�����k�Zy2�X���04��.`o1��ϭ��.�.V�t㵌W�hQ���8\S,QA�*n�3�.�)���b�+`��Y`��A���~�ҫ�G���Q��ˋH�ڧ��Nf��\pw�v�őd]Մ&Z�Uqd�^'����t�^7��¼mg�q�������������ü�l���-<�F�/n��&�{�B�Ы����Ij[�����~F�7u�T���a�d��B����`N��4��6���'�oϴ>������A冐�~�<p���w �ͼ���,��zaŹ!#u� Pc��	:��n`�?�,��6]Q��F����^x�Z,׺Y�+�E��/��N+�;4��T��B�X�T �*���􌚨G��UDp�5f�7�|Q;s�<���a������W�$F�q��7�4�@7��" �h���*:�<wa�G���۶�k���=,؂Q�}�WL�hp������a0"���y�߭�r���7A���e:�5��$�~�����*��Z���=�K����(�g^����l����wD>�x�Y��l�6�k]��B�:��α��u�7�<�VF*63Mb���n��B�m�%i��f�BEz��	���� �ls>#X� �.q�Ր�)�ul�kʴH�s���Q�A�&H0��;���=:��m�pQ:�����^?t���޷�N<V�l^�k����EXٺ��;.�o��zYwƝ�0Ư���DK&
.{R�V0������b�ܳ�N�׻�{���b��v�G�Y�B7k����9���/���^�	��ԉ���os�����0����%��Q)�vF�/��wY�&��WlXu3�}8%a����ž,�?��uŹj�*�'lN�.�U�,zKֺ}y�ݵ�?��<(v[IjRc��a�+dY���	h]m f���m�g�^��?���-�Q�uL�yBb��޹���O/�����&#|�V��=�hb�ǡaK�g�ӎ�Cay�p�O��Mg�Zb2�n���}o��69h�����P�S�lFlk�򿾕�8ϯ�8�5W��d��-�<�U�����]t����"���yȨ�^�txx|�?�c��p���Fق���ך�Sކ`�E��:0O�����j<M�u%1)�"S_<P{7�O�\������q%�aI+��<A@�0q�ҧ��W��a1|}���C^z����uB9N2����Y�əq4Y�((�54�>�B��l��l�se8���L�x��+'RZ{�		�Fp-��|��/��?\*y|�A+̅��GQ{����"���'r{%�zX�6��#x�E�c��J.���@�[���
���}0��-7��T�Yj}-A�CNg�NX��샩�%U��X���ȣ���]�[;���x$/F�BP�?-��4������v�����5�y�C�nw�kg7�0� 8\%���	�+Q�W-B*������͙�a��G��ԛ��!���=_M�h|h���lĐ�=T��Z�ج~t��sJ��D.���S�_��:<��E��wO�����uU��0b/3���+�FN*��M@�_��|4��o�����l���2ȱ��\�}�kE��	Z_�k�{;��3ӿ2F���%���Q�C�n�/ևH�!�26�{������Sù�	a��j�w�T����Pi[q����45����i���Ј𝋑Y��2;v��moo/���s	ƖT�E*��r@\^�a��kF���b�K&������{	�o��}��ct��&�g�-��1=f����וUj����y��� ��u�	y�wp �(�/9�\R�������l��ԅ��X��B��k�Z'r�8��Ki)1��e�7��+���ѯ�>vh�����Ha��ϋ���$ߧ�ׁ�K�V���r��Uч���/(~ⴇw��Ŭ�����@0z������w��k_o;�&�<8�i�����?6H.�L�_���򪱴��e���M��?�Wr�S_f��� !K�	���㙁۲�,��,���ѢơL�'����e��Z��0��|�	�(���5�F����-��j
Paܵ����r�^�x��������=�U_�������y���M���ECx_��к�]鉼ԃD�e����o��W ���[�0��Z�I4X�b�WJ���t岱��}�%m5E	/�
��m,�� ��jֺM#tG��������&J�K����� �����ɵ!/uQU+�J�Û��l���S��O�<�I>Y�O��{�छ�<��O����=X�g�7;Sl$s��Zd)z� Ia��ݢ���=ڸreE�~x�Ǝ,��$Ҡ?R��q�}���1��=?�x��6,?
0#�h�lԸ��y��
��R=���8'i�Ǔ	�W�]��7Ҧ�Lr�t�\�|���;3.���1ki�E�F���-��O��J�*O)ahe�G�\-�,�6��51��S�Ŝ���f����9�b��D����ﲔ�~j�=���^��9i��f�~���}�a��K	`���	5!�����-�{��vU�R�*H��M#w��C�i��P�)i��ςDRqh��dm�R�7��'��rOk�����o��,��o�&���3���v�Z6�B"ǔ�F��I�/>S'�����n�a��Z�q�����|��x墅�ؙqx�叠�Rh*�NQm-&���eF���6��z0*�QO��;��[�f�����o�מ
zi|�|����1lƳ���|���[Oi<�4���v�GYd��'��'�:�xc�H���݅��*�^�iS���
��:�h���9$����wdN�Jg���Z�����Bx݃��Lm8�~c��v/<���X��O ��7nUī��\��$��*���ϲL�M���b+�Du������m6�Ҋ\v�^��s#��)�45&,��8�*T0���*N6Q�k�YM4����{T�����h
��\n��pJW=5���4��C����Q�����Pi��$Gǐ�n��nD:��F7��g|�����{;�9��9�:�h<��� ��z2ֽ�����������/��z4�� �&�۲�@�$���D���]4')�0����x�Ym7=�E�
p �.����/��^������8��WSߐQB�,ꛖF�D ������zM��b��/K���;>(W���N��-��������d>1s�R���lIŐ��.9�Zo�	)AHh���h��<�	�c4�TΤ�7�7z�����)>��z���[,�npN��O"�Q���T;l4�<�c���k|���|��Q�[)��QpDI��Gţ��%b�3�y��e@/��������;;g9:�k9�D5XƝ;D��@��5oi���
���^����:�6�r�QZ�܊����L��7 ���V�V�.�&]�{J�s�2$��ʊQ�n��8Q����ߗ��=���F���/%���Zjyw(h�p�PV� tƙ:�p-V��o�� �"t{�k՜��ly���T�n��y '�R���u��!�I��.��d@��hY;������ew��T��ڏ��
��Ga���������{4�I��׊Ȧ�}�(

hi�%�o��N�6q��ݻd��G����2��/�'�^K~�"E��LU�� _j|�X����$�<��K��߻S���6cUa;2�4�#��{~�$�Y�?B6��v�G˅���^h���!����7�&D���"�_qYK�}B�ҟ8Ű��I$Y�z3�W���~�1��4��	�$�M%���e>���8����{Kfw�LR��������ߝ_;��Sk�����'��ӳk'�1WlLQ��l��`"�O��m���RHY\Γ���ۼDZZ�9U�[�Tz��p:WO��ܸ]�<��7]N;?�����GA����x���(������H�y��Sx��nw�S�Ŏۈ�p!�C4I�(��q���Ɵ�	P��.� d�$1����B�����^j3�	��9K	Q��<�=:X��ځ����������.���֪]V�cum�ϋjG����Z-ٮ����Ӷ;�P�PiP�<S6"ȣ��(0J1Sˋ�=.Dpn�譡l�>ja���3��m2�dJnL�[h��G�yӯ0u����x�,H_�ҭ��;����x�);W^
�T:�H��~��%�~�U��.�h��Y���ɍ8�|���%_h�P0��a�Ƹ3��!�Ci��b��ۜ��.1��@�����4�]R*�o��$�H�T����p��*o�x�)��}`7�������㾵��6u����@���j\����d׏C��QZ�n�/VO�ev�t�h�b� �w�I�9����+����:�j�*�Ep@��4��N�	�7RL[�z��x���)��FQ�č�8�|�P��S,D��m��m���q��ɥ���䢞�X[���� @�mB:}��[���y���N.�/���P�����3���'v�qye�����щ%h��V00�Zu���g���_kC�̱���
��{ ��������n�����'��g]�M\[����O7J�CI�nF1;�rQ�U?��9�S�������4q�����^��B��dyy?S���G�t2�:(�	�+�[꘣�+7�FtfgHri��j��]m�[ I)��9>���aJ8�����B�b��@�
$�G*r��L�ˌJ��S����}?�0����sc퀧�ߣt� ["�L8Ե�`c� v�.�H��@6�5��m��v�}�����y&�8�d�}*S�=�7�1+7�2�p��?u�=��V������1����\���P7�RHvo�+I)��~%�|؅�M�%;M�Oqnɬ�}36g��׳�����a��+�ԫQal��a���$b �9ݻ���6�
�3bn��\��:�G}�m,�u��܏)L��bQph9����y��4�
����AR��yR�b�O�\���,���6�իv\�r�=�=y�/N��f$�z�]D۝U����D_�����sZ��E�M����0ϡFg�N�#�����ԏ�[��$��,���1���?*��U%��>���e2��7�����S>�6\n''|�c�l�A��z���w>�x�{6�s�dax#��V	� �����M?��FyQC*1 tb�Պl���h�<6Jz�im�񑟷y��%
��؍q��H֌�����Oٛ�vE)�6��"�\5 G����y�T�1�/9���J�2�!7�}���2��Ä&�qU�΀,��&IdT`�����Q9~�xXZ^'���ީJ��R�25MX,͎��1�:�c��~%�995��°���Li.�F���{���Tp|ݪXc�7�,8b�b�Ѕ�UȤ.�s5�!b0S�� Y�w�<2af���)�HPET9sP�5�7m~(o6�K�@�m�#Bû|*�RIQt�<)�|�Q�:P[�A�3C0�&~й��?�>��͵����U�%��w�f�i����-Q���<�=Be�{�_����:Z�m�*N�{F�����V�&*�/{Ѯp��)��M������ٺ~-g�����[�V�ǿ�� ��ڟ:��w���DU�ǻ�ǗY~b�.vr� ��	915[P��Ɨ۽R�Ao�I_�-�t�sQ��O�*o��������D��16ܶovVôԤ��Qy�%bN�8���y!غ[���ѽ��I�+���.9�_������qE�rA����?3�j<~�3DAe^zڳ��-|�W@�(YR��xu$Ő�"���.�z��[0!/t#lc_��F6
�2���r�~}��t��P_�ZB�r���s>��j?��c��WtD�
 �G��Y��peN��ii)�PA ��&�[�p���T�M�
�Q��^s��}`��H%�d���f|��F�:�ܩO�T�e��ٶm�N�h�.�F���v<��ll�V�k'ӭhDf�Z1P�aZtX�	���ǝX�'Ϣ�KQ�f����0Ƨ�ُX��ߩ��}�w���ƺ��!:�t	"��2�Zw�G�=~X�ܜ��j-��{wQ��Ȇ�"��תj�ܞ��|cm�9�Zz4���!��i����[AIH�Ц&2� dD�n�U�_̪�Irg&�3�H�Q�)f�=��?�L�̟��6��
���ȤDϞ �����8����Pp�N��T�椧w��d,�;B[g�s��#�5���V^�� �K]G����r������#�o�Qj�.y3�N���w�鐹z��S�� aV�R�_���b>�eG��������Ʀ�Zo��D���Z_�Hmb�k�39�[��Uv[�����

�K�&$��?ݭj�K��3z�����4sXUh��a�����-�k!J-��zQg��k1�p��`Y�ͰM|$at����XH� {g��%r�h{��FX�C����}����h�`�L���IJ���WJ�
M)��7s��̿[Z,���}�-1yg���S}��g�0 /�H�*�R�RȍH��'�ZU�9# ����X��'�b�ym�NA+�P�)���`��?�zh?���{��8�����Lwq��6�O��$n~X���|\[Ӕkn��=4�?$�\� 8iE�шY��ƄtcB��}6����%�����Xi�L�D�0�3�M�D/ϼ�F�-��f����b��.�7�\�

�N���3��&�D� �D����HBq�B/��S����3W�����+�s�}�]L����*B���Y�o���w���:E���Rk����l-B��O8H��H��Jpv�y=�&��S!��"*)��':��2����kW��	2p������c�[��m�yS��r��Iu�GO2�VC�h{K��Pip�p�t�J]ڱ����vr߼
�1{s�@�X�ԡ�����#��)�3d~s�B[9ݎb..�L&�<j�|؉0O�۫:#��Ol;Hx���(���j�_�ڪ�8��U�̃K:N����h�B�~uy0���w�nG��E�U���_����l'��(�X" �ұ ��k{�q���}�U�ᩛ��SSS��<����@i�:���μA��G��<E�ؘ/�sM"�����Tr-�i'L��?�'4��R�3�y�.���a�_y���6���&��JR�h��� gb�\����-:-���V��������r��eZ�#���0oT9��#�����ѵ[X �o�_|F9!a���|����<{��xĖ��䊹�����;@�@�LJ*��.�6Ń�)5b.o�-_�=���W�״�i�x:713e��Sѥ�X�5�s��1~�\R����5���n��E)4^o���;�c�:ZL.���r�ςikk�Ꭹ��i���V�c����trt�ˡ#����lua=�����%�"r�x��\Ѭ����u1����e-9��Cm��(侲e9�ޚ��O���4��<܎��@_�����k�#!;#ؘ�o%�^@�*��]&��KO<��8qi"'UY�zS>�d�u�la�_�����<8���׶v�x
	tM3�+(I�;sѶ�)Ô���P�@���{�]�(gYk����h�	dſ|�O�|g|I��s�����:06_'�_5Dqs�d<G������ʗtB��ۯ�Bt�̄s����.���,��͆'=$��Cj븗��b?�Ln�u�{�|�2��b�m���$���;85ϩ��'���PM��L5��I��?Ύv_K�w�m�]�7������#n}=e��p������6�"�F\���B#�"C���^��!K�SK��Pf�"�%7A��Mt��
�n���1���ƶv�=!Ƹ
��c7�W�X�yq.��M����Ìٯ}��3����i���Ѣ�z�XBؽ��|�?�������lA)��(I����vS(H�e�J�rL�y}>q7�VJ�-��1^�
G�-���V:,����
�iqs���|ԑ5��da9g)_��.#b{��4=��������{�	��6�ȅ�����D���(�3�"������223&�4�@HS�2�����Bv�M]Cչ	��Djs2�Z�s�]�Q9�j�9vFT	�<X�Ŷ�����0���c,S�A��T���72U�Oa^p'Ml:��������*�����Dp��pI�"i6�)e���@��˯���&��8�p4�^]5���xo�F���tp���\?|r���D���V�s}K����z�GP����~Ҝ�(��=��5���Z����<��/��g ���I6��h�s���כ�6ܲ�o�ݯ����qT>���C+�u%Y9���)�Q˛��=5u���E"���[P�_҄;52��F��>�:��!c <��*����hLK�>QE������;��y��W+~�
��O.<c�ݏ�wj�n-��{(����^ݷf��'c�ZBQ�T@���r{%m撥�MՓ��ذ�ھ�#��y.j�C��5�vA�b$���m~$�4K�T�>X@U��N��d��w�}n)��{��/�>���.��*%/$7y�)�{֛��#�D�r|�K���I����5݋�9�.qp� �է@�KzO�>-I�ܠ&�H����S�y�ܰ��!"@7_/�MMO���oPe-�]!0mZ��ir�6"3��X4�#/�AU�v��l�&PF�=}�9�=b��~�ϙ���LM.��ۣG��##�5�Տ�,T�� rh�)X���p�����5s���\�÷F�
;:���Q��2ܬ�열��~,� �v:g����\�>�ᠷ:��V/�O�p��"�yil�X�Y��Di�~�\�j6���&�R�Oyi������m!v�]�*;���0�Kq� P���[n��EV�Sc��b�ge��V�`1�r�	љ^V$K���#��f?�7`p�cI}��[:S(�%���1G!�D��%����j�����綧��Oq�H���1��m��~����Rh��d���p�{��Q�7��7��n�c�o�wdJ��Rmh�w3^�:�:���jF����)����P޶-7��P٣0��#踀���z�$���P��-f����\O�G0�#��JYA����]h���f�S7�Hi|���Y�>\�p�-N�����b�ddأ�d����2�A��:��/��vM^	>�Rj�b��Ge�e��u;m_���;�`�*�@�[<��3%�]Y)4N.����uz�#����ww=�XRKl~��6�q};��k���.��y�[���ΑG�=�7z}�=	�E��;w�CXd�r ]$����W�T���E˺3��}}�Ȇ$��n��Zͫ5Z����t��,�=#��sMaX�>drZ��~E��jp*j��
�Зu~6h�߷�[;�%&!y���QB�-�ɫ'8P����M�ҝe&U��MR[:���
�b�5����*QbO.`I~{�t�bY:�na�ǘ{�]}���J�U{��M�- 1R2����G��_�jA?���X��U��t`Wbh�v�S@��҃է�����nՒ'oH���nv�}w� &���g'r`��x��z�eN��}~�^�\?<Oq� �#���bgM�AAv��6s���I���]�'x�������R��!�(�W�*�"]�	S��8�~K�%��5y�GAMT��s�(f���͎�ܦ):���9�{���~�׮���[�G0s��G[%G[%�����់l��,�iYqW�+�p�#�g�1%��y�`�P$P�d�s�ģ�Wn��4-$��^�	4bE�>\b>�U��/�Mhhg[A:�o��0���hWz[�����*��9w�]���]������VÆ�Rj;Se���(�Lz��?���҉d�/8��(�&�j`�~`΋+����rnG�u���}���~衃i�>`X`��m6<��;���N��h�MmZ~�����Υ�h()O�]y3�rVo�p�C�	b�>I�z.f@=���ԩ���t2ep�*̐7ò�K��h�R+�\��[�ݝ���%��b�Ä�y������=����~�ط�����.!�C|���r\�x���zp�72`6���/~I6rJ�������&�i}����)��:�C�Qs�W��[I+�7�`�_1��A�?رJrn��.�{Zr���<����Hc�D���׻7�cUĝ	ɳ��͍�*0����w�U����rm=o�8���?���~s��,����}�;�W�6�s-�'�.A��!l��m�s�y�ؗ�L�7�l�\I�ѝ,w�kF�`o��mh��Ѷ5,R�x�D�wi���m�Z�=b�#6�v��j ����{k���$e���k��kV������B��ŁNL<��+$���D����1qWK3�V�,�L8�߅(��m�(�/`�IZ�P�ƙ����̒��I����8��v}Ӂ-�*��
8�9�٪�{"����nU�w�2ЍC<4GD�(���J�i��j��<J��o��ٙ5�@��.c4�_���v,x�~�����ۙ��R�����鹺�	�����	�tAH�P<I�u c!Z���D"�LYQhH����I��@+RZ2V��z���J�����蝚�ob�-w�T��8O�y���|��=a���͹��?��d?� �М�<({��F�_`��u���#��(�V��g-%�z������j�y�-�;
2Z�p�M������a^Ͼ���T:�3�����r;_���':�U��"iW�+N�ΉA��lƚƨ	�z� @M��Q����81h���_�ܣ
��y�Ϋ��1�`�>�� %q�Ƙ�����p���d�a˭�K��Ki�7ۣ�&=�5�jƒ�d	��wzS�����	�?Yv����z�E�f���0G�[x�H3���}���q�+��Zq�	U�*C���f<�{S�3�au�&�l&�⇒`/'�@�:���q�A���|�K	�H�D=4J���^PT�Y`��D�O���{}���of�Aj��*ڇb�ڹ<��������Gҝ��U�:��@�>������FLە���V�d����8��GKf6�5���<F5� eBN��;{rW s���4x&~/F�)b*N|���M���p� ?g�o�F���糮�J1ny��ȕ
�K�h4J��n}Hm��:��2���S^ac�!�{q�B��#��,;so�'Q� ���5B����`��/���������6��|#���2�՜
�;o
���|�[��xF���К��A:?�EI�������)�q��ũ���$W�~Ŭ���̐R.�$�:~�p~�\שa-N�[�7���;
�U���w�pU�O�7�H*`��9��Z�a#�v��D�6,u�v�i�f��y����y�[U�yUr����y�_��?�VɆ�Θw�]l4�0#�12|ii���k�l�p�!h�)a�m�^
tB#�Z搪�1��X'M���;ݘ���0����˞P�<X�Q;4G9������ N5�h̽�q�R�;Wr��~wT²����̅��q.�f5����b7��-O�)�x_�iMn�zA}��@�Hr����r�*c�3����f��sH��`�2(w��9�������;��ђa�f��u���F��<y��O�K���)�۴JW;�D�|}c.7�M�rn{�b8��,��x����;qI�?;U�&����l�H��MUu�<�E��Z�X�'<����	��I��Z�Y'�r��KmGA��f��8�|^�N��I�0a�Vޤ������u��3�7�P�'����yX}l?���g��[��X��}�t��b�����V�~"�P�AD�V�^N/�Y�(��;�ABۀ�'N�'*�oP�N:pT�W+	���sK�q*���D���Ò��1	��Z��@����ӡ4>ʔz��/
�^���k����|C��nM��8�7����N��?sZ�5����S77�:)#uw"�*�`wڼ�gb�tF}�b৤�Ů)W�Hf�f������.oy����sH�ٕ���*��DI�bRk�@(i\��^DZ�D#r���(_s�f�8Y�:WY�y���qi��A���/��'�6�s�QM!�3�A�vP�W}�AUN��MF���ت_�pQ%�+����|M��M�7��XVU��[)<"����BK�f�G���Ό�Y��w7��y=�5�=˨�p�P��P�|OuyЁ�m������-EW����&���z��9����9HpAV����a�aDޕG��:.s����TJ�ރ��c���Ԙ����� փG����h ���xKZ�.���s�qO�Ϲ�fN]7�#��R��@�J)�s�����:�qh
��:�������\��\�O5E��S2e9:cZ�������	U#h���3Q���T��A����A]�|������#��ű�bf�n������bI _��41���}V�� �_��>v}�K}�6��;kO8{|gDnp�q���Z!E\U͞3�uU��ϙh��)��@i��% A	q/���t��U]7"�#d.%�6Sn��VL1���0D9(m�$CR��s���?��l�u,N��m�=뺈�I���E����/���W�?��|$~�\f�k~va��Q��E
��(�JT����]�&�n�3�9��(#$1��
i�eH��Ǔ�n�v�9�5l���&W��|]0)���n�N>Zo���[lzZ%�./',>$�.F�׬������ߔ�&����s]��ư��tƀ\5�9�P�DK��i�V���R��\.筎M�kX�EV���&$��~3�B~,N�I�~©/�:c�1�6�h"�I�'vU����g��o����x@��tD�*�1I�a��w��R���UE�W*�I�X>Xn��M��PW�N�i�5�<BH�����ߋ�5�6�Ct�U�b'+	e=��d��eB5�,Ӭ�BڈUR��9�}gˇ��
^��`�d��l?��}�\�1�#���Al�q`�/�N�3���Ģ��6�8y@%�@����m#g��Cc��%�����˷������`Y/JI(�Q�f>6��	��͸Uc�\B�\�~p���|x�+���������D�S�(����k
�E�s~�������ZBCS9�@�K;�`���!�Q�_ID&���$n�4�
ۑ�`Ẃ׉��+6�d�͵%��7M���S���� o$?�EC�<�u���N�v�j<o
�V!�t��O�𑆰���Q�>�y.&71)Ϥ�BU!���=.u-�D��Jo������]� ���ݫe�M�;YI����h�܀�>�lZ�;���X�6c̈���f����yxr��aD$P�z�ʊ��&n���� ��*��Kf������/kA��~��j\�D��^���{���ԌwX�I�\��rF ,�:|��!�1Rٙ����~��Ap���o#�tڲ������߰U?��'����Y^�qI�P���'�2�	`���Ғ>�J*�F��-9�2j�dU��f3=�@t֍9�Ŵ�<�y$�p��jӖ�ܵ\��^g3Y|7B���i_���xJ��h�6����^P���iw�1@�Zs�d���P�͹�G�w��{H�9ʶ����%�M1���_���?�*n�o|� ��,/v�˯��r��\�qU3i5+�5ńo�[*��V�����������-	��)N���#��Ž�n�D��.f��z�<������ϔdIm�a�܄޴O��쫤����o�4qG�Q�J�P&erV��	ei`�&z���M֟9��I��(���f��Hdu�}[�0ź���>4Z%z�l�$bg��gjs@��Y-��ר�g�B	�^o���7.pO�4����@!ta�3�MSj��1�5��j�]�V<2k��:Ǥ��j�?ЌݐK�d.#%���m̃L#:ڕ������[�Iob��{��uP"�[;:~ �%lR��mtq4v^qл�-.a�Tn���d�5e{u�6v��
���|�g�z���\�i����S������ʣ�p���vr�$+wzr��p������r��WM�Y��]~M�-!ǐl���%�?(n�}&#l&���`!D��$�W��S��L��ލ���z���#�,�
<�M{���1�*�p�׏��s���i2<�M�j.�Պ��d�.<����K�̉�nY�Y@�4�BrTת�j�y�1�`ǣ�>�s�D,ICȶ�ф�
���|؆��߈���=Oڏ�]��ZE�K��j%��(~UA:H?94��p��0�We�&�8^�q�֮��� �Q`���%�T�U�$��rt\� ��������ee��]�c��*?˷��*ꎪ�H|
5ܭ�� �oѧ�'u��-�[��N��?p��?6��/��o�~���oG
���6������>׿9�#Pߐ� �Z3��ꥮ-
�Yݟp�@��6��-�/���y���zˏB����%I¹S�Qk��9R1Pp�x('���d{p��N ���=|�[p��l)/ے��K�r�I�{�X�m�H��[��ɼ=�P�M�<�����h����4RQ�\����SE��-'����7�tl �:VCx���s�0�o4���~Q�+.�(�u�h���+��2/����eP�7zʤ���:�y�C�x�ɾ��al�[�^q$>�+�$��ƳԎb�}Wo��^�&�#,yL7�|Q��1��>'�R���&��/d-��e��ݞS���;��ށ��Լ?�K�^p��Up��ņ���AՉFآ�L��7ZU�,�������=WU�&p)ɜ�p�	�V���cH>P2m�>�^{�P��.�}�{%�M��{ji?������tUx�]� ���	��:7��!��jIT=��0,[}��>�W|:L����1�)�˽%� Jx('ח@GI½������Z$���͛ܜJ��<JY�Π/º����@��ӑ� %�����Q�G]a�B��R�C���&��"�咑F�����딮kT_���D(��=��H~FE��� �5�5�lt&K�M��j��]=��M4��$�N<v��^�)����LG4�	��]5K���m��d�~��:�;D���u�W�Qȍ� 1=��xL\'��e�j>F3��|�&�Ξ����xm���(����H�'����*��v[N�X,���7����C��T{������T2ސ���D_D�ꃁ܏��}?|�6�M±��~�X��i�Y]يԂ�=��FN�]���s��R��R}B3��^�'�eJ=��n�����2��_Q[���S8�֓�%_H�{M��o%�2tAa�F�^�rP6c��h��> ��������7f��p�-�Hxc|�/Sb̢f>�|r�����:���x�|!��cK�]R��d�_KD�)K��r���/P���zGߓs�؄��ȇ݊l� �҄���@�çU�V��&e~�*Nk�3��ӝl�(�O�A����~��7>���~k�_���&����	��GX��1��-��Ĩ��R�F���O�I7k���)�ږV)'�evt1�{zi�Q<�{!VX�P�ӥ�J��{������iF���O���!�+���V�6tRh���P�!}Jo�8pr)��=�R��Fה����F=���j��5B�t*��|k~�-��-�\=%I�T�"B��'�s��wG�C������۳�.M]�n"���W� �dC�ħ6��͇}��W��\���+�,�lH�����d�v���|"ؒ���Ʃ��n'��*!������Mc�Kzѩ�"eҜ	!Z�KT�{<R|wWf�J�����@��{P��ygCХ�R�>��#���}�lA��l���p"G�;|���W��Ŋ�Q�[W���v��)�ݯ�L)�5��v��gB��d��]y�t���P(4n�\o�8�I��W�|� �9�������p ثӕ�{(87������d�2���.+�0Kq�)�r�|\]r�M}␘vH��q�[��&�"晐�SFq�>�/U)��@W��f?�H�H����(^l���T.{�S+�8K`���b��pr^�dW�lQ;�::<U�?�^ihH�<�@���0�U���R^�bB��M��v�=*^���'���Y�7������� ӭ�6����'G������_$�s��*�v�vs#+�iHm�����a7�X+��2E��-�P�[�����g�����-��e� ����=K����:c�V��r�͔���i���"�A�,۞n�]�f��X����uhd�{�[�#k�2�zD|�4��_�h"��YD˯��9B9]�(�.r�J�{÷6Mg��+�:Yo���3=��z�N��$��2s�0B'O�9[��������%ȁ����*�覦T�̳�?9~�l&�C�0}%Y�C�_��e��<���qgn�δ�O�W�q[oV�$|�1܎��l�H�pa*1^�.}'�&f9�l�eM���
�R^4ԏ�U�.m�3��˫&a�?��Ix�*<��FX�����d�a�.Ȓ;�\�N*�+},0�JGC `{�u�2
gt�[��	��Z��+�T������[����&��@7A;���<P,P�3�ٞ��U=M2� ;V�B�	EK;���n�V��+�C�J;�Y�0� ���$w��"4��g���R����/-Mb�z*������/}Te|ޒr��pVw`"��H��@�%�Z�W����"�Zuז��aOY�:�9u�J��ih(b3��jo���E�ڽm�J
�o���e���b�d�'U�4t���:�U~D�I#�<��MjG��������A�~#-D:(�L�ԾW��ۿn�k�dy��X�j���;EQ�P��/��U�ē�6vŚ��a�^(����)�
�%��A�zm��q�)}�3bF<r��y�9*�����W�6�M��߆$.�*�k_"��"1�MeH8AcOy�BQ�FF�����|�3�bh?`�-[Ce��� ̎T؜˵��Vy��$X��;���3ᇗ�-6�Yw��2�ѓ*�����>�:��)�^	��bs��)4����<uOG8�������/���v�h2�M5��&��7�N��S)l��4�{m���ԣ���]觖3j�� ��s����/���@C�����2�(��n���BC�_[/�M����Z�J��in*% �+�'
��̪'��q{W��,�J~ji:_4zR۟�Jͽ�m�Z��X�QW��JҖ9��d/�u7��u���hj�P�D�l��Iv!$����T����E]̸��/�����2�#�^m2o�?U�q����Zn��=z.���*dODW���;hZ�&�S�H^8?ޔw�-z�$��I�._-/����	<[��'��<�c�e1 ���ͥ0+���<`��0ܖ�U9���б�Ƌ� ���CA�Ï~`��\�f��P �w�'1������ڙ'���w��|�۷���S�A�Φ��|U�e%a2]������hB�w����0����ҹ�^4�*=!��|v�8�k]V$��3��W�$��w9I�x��D�&L�Cl�T갯%e@R�+�����C���y�n�ԌO�h5�s�扶ӳB5�d%3$��8;��M��;�=�x\�+;QR���-�ܜ/˜_�a��\���d�b���%Yo��Qb�q7�Ia䨰Ƅ/N��t6*y���}%8��S�<M][[��&�<�/�Yr.���t4,��uS�>%d�~x����ji��@��������{���՛t�&�C�Ŝ#j��m��h����;�~����'�^\�ݲ&���o��-2C��2�I�Yg�hn����]D��@T�Mp1>��}��#��OĩW%���e*޹���]m�+���T&v@�^0/���]ﲬ��ut�[hN<H㇉��Сd�>�%�՛��i#�_<+ /����Y����B�n�[������}���sz=\�W:ϓy5�$�%��U8���%��Ť������U���k�(��j�ݿ��E���Z���HU�j`�����:|# =5.x��B��.��Sy����l�z��H`�#��b=��x��"DQ��#�Z��s���������8y���[<4>R>��VF0�<Q ws���M�ο��;��k�~���7M�7��T���kΫ���w<����:2�E䧼�h������p����Hź#9��`�vO��P��+�i����p?b��(�`�Em���n(Ky���\�u��ݬ����a� pD�	�՚��'���K��� �}%��r٩:s��e�9��*��9y٣C`<$����*)`n���6i��c��gc�:���_Ȏ��JP%6����[o̗��z����'Z�<(�P���Up��U-�h,�t2�[�~��!�7�Oq��M
���#�@��N�k@}��9�X���
���k�y8�AJ�ʙ՟��óю8���\�}���L]>a{l��^��n����d����Fz`/��ma9��4�?6��A�X�f�B�y�B)��WU,�E����P��6q��|�~_�f�����m�Z��A�Py$�����8˯,*}� :��Yk=J��ҍ��g�����56?׮+�P�����	�~�AȄ��@$]`	���P������-����{"��?�G�i�����Y��ʉ��>JxW[�c�#z�+R�]Ft��\�ͯj��|ZU+ːoO��'*b��}�3������5d�����+���^
�d6cTܪ�8ּ
(,`�		럯� F@Ԫ�,H��hmE���ߺ)#��a+�ǭ�\KZ急�l�����ߏ<��l�M��tՋv��ti�d�(J5��g����t��oy�2��[���^Nh�n��w�>��{�i��+�rDժj��q���j�7t��7�b��-�c�ڧ~
dWV[�_/���sa�����y�ގ� )Q{��*k��q�H�n]s��-R���-��D�x_4�����%��o�t�NS�������`o���;��U �>z,I�J*?�Y�G�W�i�zኺk����Xp�*_C�����b�����	���*��K7"7��f{F��^bI��UI� ��\��S�׍A!�ԉ�!� #GD`�5}�w�L׬ڣ�sy3��� =��o���a���,Io��[� �҉�_A�������T�#�'���z����Aav����SVlM�z��� ^yϿ5��D�V��D�I}?��K����oDu�=ءd����r$�\� 59�(߶T*J��fO��W.�
J��.t҅���У$�1��_����<n��~EC�4��FQ�W=�pzz��j̺>��nK�U!��%��Y�Ω��8�%���˚;l�\�T�>U��H
uÇ���#���É�^?~�y[Ki�WA��Pw�i����f�t C����lF�x�ߞ���h�O�՝���Uo��u�V(Rܡ���C���ŭXq�]�;w�����z��ߝ�g2������k��J�׈r�|{�"��쏞��o��/S�Ѿ�䛊��X���U����A�Po��Y���5H��2%V��3z�B$�l)�����I��;����k��j5�iS�Ǵ�.�ji�j9��▰W�o�:Yk�W:֥n�:X��H;�B�ۈEz���E��&�k5}ҕ"�H<#;��(a�����ޖ�&�D8�6G��9;|_�f�k�_��kS7@$�T k�Hv���t�`�8��w�]�:7쮁a�[����J����\m��r'O�w.�k�Ȩ�P�xՅ�ޫ�����Cwl�~�� m$x�����BHf�e�����:րi��qO����Oz����њq喾�=}���R���5r��#�8�^��e֪��S�Y`�1=��	yeeZZ�9ƹqM�4u��[0�K|�����(��[�<]�(���I�M�G���ѿS�����^�【�g����Ɗ3�Q���]��ߦ7�7��g��l�D-�-��1� t.Z',��2��Պf���/a��ǰ���N9�"4P-��3j�l�v��﷗�j�5�:дE@�Q�?4P_Rx<�>v�����BƸ��L�c�)=x4�$��H�[#����
�g�l���)� �/��{x�Ң;�-Io��q���ז{��v��f�g���1�[��	,�b�@�y����p�E�GR�uV��z|v�ldg�����w�6��P�u��Ϲ�����Zk����ǐ5i��q�=j�^/p��	i>_
���a'�ka��߮aM�?��>�+��d��R��`鮪��6g�;������Xp���|HCwU����c��Lq�ٯ�O�ܛ�6����Չ�T�Ld�YMn��Wޘ�q��r����_��%���<���"hwp��Q�(��BO�_̌}��makh���QTU�c��*T�<������&����LS�KmP<C���=..G���ݮI��L��acC��a�L��f�e�H��XoO[����Ewi����a��~�y �R^��.��b3^��u��@=���_��߆�@��3G�x�)C�d�;<�67�`�����ef[I��6_�X�8��?̖��/���v���.���i�FV�1�0���H�p#D���'xP$�e~s� Yش^���ϻ��_�:����]�1���D�+dx��]����rU3����A%}`��F�u�ju]2P�1�V�ߩX�4�@����������ҝtg�c�,+��N��A�JQ�Z�*�["���u���JUe�;�-#e��-����O����ڭ[H�I81 �,>}nEX#	D�����g��ae���o��Cr*�i�U�~`:���Ӑ1K��hRn�Ms���/�/v�8��,V_t۾"�f���Q�C5Eee�'K�q�h~��7aR�}[�E��#(SUA����5��;����I��UQ�qX1����y�I9�1����[���-~�{�!���7{G�`�1r�^��eD��Ɨf���e�}�J���ʍ�~ͬ�Y�G�o�:-���Ս��6u�lB����3��\1�*sЕ[�-*�����[����_w9��q�{V��^]�xrgC���?p/I�4�Y�����'�,Ci\S�>�%�~���+8q���F���#��#}��so��NH��9O[pD�ƭb㔛��El�(Q�ߜ��f_�)ů-̃3�UȪ916�k�\w@55�/ŪX%�/�L�a�tU.gzx��R7�dɞ',xzl�m_�I��s;���b���U|�[d[�'�6������*8i�:��%�~?�)0l��c�Kog�E5�3i���":�ٴ�d�"�m�ڄ�<ԍc���I�ros��j(6��$���z�����1wl�~��a�j��%l� j�y�m>؏�*2�'�[��~&i��h��y�@��Sӝ~�h���>�W�<�����M[(0�g5�=���6���BX��(ٷ���	�^�o�����I��6I��B϶���T�������vg���,+�,f�����U��y�`Iu��5���c	9�	�nݴ���(��q��M���x�ϙ�u����>`B� ����mUa���_-_xr&��)��eD�S��[&>
����|[��^0Ll�Kh��u�!��k���f玜���(3�q'o!F��Ʒ�'�c��_�t�UK)̙����C����|�»W(�B��u3��V >�	�8d�{	.�U�,Tj���y~��g4�~DJ��'�aȵd�E�N`*v]&ᔙ9�,��U͔g���2'��8�|C�gR׶������ LY2��v��X�N@@Pm9G�y9D�nL�+	S+�T{0.�E�~ ����2ôy=����D^'V`����.C)р���Yy�ƴ��H�T�H��-:=�nɌ�n]a/�X$B'~K��d��@N�cϪP�_���z����#�߁C,�XϷ����zneIFb�1����7�����}#��I ��i�'�*��U��!a���u��f������ij��mhZ���7��yI��dx�&."t$�H�H�� Բ�9�m�7�,�k�TL
]!��)�F:R
Y�2�9�B�/�����+�u���Aqyy_$�:t�#��_�+���ő��r�LUm������L�	��p����Svpȟ=�SH!b�GD*�[�|#���ض/����\Xx淳Cw�ϿYƃ��u߳�����W\tp�))�5�>���;m�-�W��6�zC���y�_����0����N�Vs�>c����AFH�!��9��Cy�x�������ۢ�WT׋��@�Z���h�vaF�W�?Zo�ݮ~�Yj��.��8���"7]c_�k��V�=!�>!�o@<j�9�آ�1F#���c�x�����8�f�8�ư7�GQ�G����� ��Tr��q����x/F�8t��Vy���*��k�;Nz����w�p��\bfcM�Sko�U��n�V7����J�jVv�pt�?�)ָD���n�\�o\/-���:+j�N-��J5��w)�:��L�W�-���I�,:��k�e�Qi��c�6�K`
�΅�b/g����UA���Qwy����C�d�^i��~-L�t�nX�H�T>��3~p�.�_b�mŸ@"d��п�Nwx$���5�����ǃQIP�������=�of{f���@a��RR���b��c#�\� � Qj�X�	Lt��o�LI��!�N�ZTy�]�s#�'zpQ��'����Ᏹ�[v������[�ܟ����?T��l5Z���'|��Ϯ��ȴGH<�߫W�E&&�L��ftv�i��*�F`:QC?�X��i�Iۯ���J� [jZ��y����VUw��� l�r���8�c��͆6�<�8"tы������̋�:���ҒB��쾔��1��쯟�|#~_�O�����8zGB��~u ���,��N�<oH��fk�|j�3��a{��ß|xu2�� �U��.���[�
���J�8�~�|�C?c����z],&:��_���?Egyi�շ�HS�c�QclW��y���4��Ђ�O�s�Ǐ�_�ҫ � ����`��	]�#�+�*�h��Oc�V-������ m1���5��ZӦ�<,��m`��r}t4�/<.�W��õBN���T��T�����d���:���F�蟧�'OHl1*QH����\h�Oa��U�����Bv&6���Q���q���(�2���@}���Ϩ��w�ͫ���x�끫��:��8Z��������Iw�/A鍺���,��X�L-�!J7A�t��p����1�1���E!ť��,�a�M����h�� aJcJB�Ll:u���5���Z���@̖�9�A�Z��Vq6>\�ff�v8St%]A��}X�k��78$�2�Q`*H� �n#&X�̹����O:��&���,��Qeyb(��ě��N�ھy'w��Fd�J�HOYy���_]���`O__�7�7���?�ؔcV��~'���6]$Wգ/+1#���Y���N�YII6�bΎT��������caa�����T�j�|VU���{��>��e��5�ڧ��}6�##uV 41{�0abW��������� �rE�()ޱ���1��{�����T�������v둈����@���rE�#�m��Λ�pm�qsjb�p����̡�`gb@P�DA� ���*k��E���vo�	=���Z_������"4m����Y�:&��i��|�m�%}�*�a�$�;��_1��ly����)���5Asȣ���臒�(	��e=��D��'@{@���N��m�A�O�]g2��[�T�m�`'�Ev^۶o�D�M��l<��Mf�ps+\��T�u��ؖ팊�rlD�^�;�"H�:�#ۈI�3F��)���rJ@�O+Z{D�������O;|��y������/zM(��֯�0��$(V�7}��h�ЫW̦���D���>���̪��Z7qW���H�Z�(ԁ�MN���㡡�X3K70�݇��������
�t͇���r-Dy�'FH�1��Șa;�[F
��ó�{5�xM/�"��:��a�tv��r�]�-
�#�q-#|��
��F�Β�\���*j7�=r�G�$!E��C�i��Lp�Ӡ�	h�[s�+ ���֢Lh�8Q��A���(G���Ä�G��R��,$;����3v|V{#_Y0�t;�-ꟃj�=��V������Տ�>��(��$1����!M��2r���i��MC>���\�Ș�<}R�-)�˶�P_�Z��	&�^,n���>��H7�I�p����:�j�Ս��������%�;�H
�̱GCJ�\M����1�����YQr!�߽MyY|�{��)�0���� ������C̱-'�JH��B�"׷e�v�FPL����(}�:%A�R"�_n���5T7���	�{�J�VH`��ǎ�`�.YNg�Hlo�j�)�b��5��w����@�w���S( ��kA�Ί�Ts����x��8�P��v찵l�� ����gO�I_ǈg�:(�Y �[���������`lO��<.3��76��9D�5���Y�����V=���_�|��n+v�.���Ș�~)U����g�5o�J}�"%ƻ�z%#��?Q�D�6���8 �U߇l���(��_H_�sW4��vfr �bE����2��Y�0:�=j|�R:�'sPs������nL����"�G6%�_U���@	!��3�M.-�;|?�����.�w+?I��N�*|�j:�q�0�2}W6�>�x��@vGvf~Rh��Q�����,1��`!b,[ws�R�W���w_vW4�r8��'���|��HUZ?�q��G8���������C|$"Bh�g�˓�Ƨ�eN_.�<�Ľ�%�#�t�^���]�c!fh�B��-d�~g�|�m�!� F����jϖ�"���~���Q
��[F��l��}����;��ng�ʐ��x!�6��s��(���@@�{dz�F�D�Xp8�CU�F��kd4_����9����U�ݓ���U٬�>���ɏf���k��o���%`����/�!���G�b�p�m�+#���{����!�8I��-ɤ�=�&sL2$5&*;��2�rdf9@��s
��Lo"P~W�J99�Q%�x:�s�O^��_ڳ���9|9��D����_��<�6�9D�u}�����*��	��vMpH�ϵ��J�b��m���7H��9�
���|��;eF�.��=c-�z�=�~\��a�E=��5�6p�,�ujz��X9dEl@�	֪mE�bj(ƶn��d��T��Lw?���	�j��/�A��@�[s������8|��?�K=�0��!+P�c�#�?Q���7�}�G��e|&_�\.k�ި'�Q41�tnmi�%�X�׺ :>�~g:ml�/;C��mD1M�`��O7��l����
f�^(q�2�~=��8�-3�;��d}V\П����t��Y)~ƿ;�4��~Mm����d��Ζ ������($2�w��{s��XMt���\������$pV�d��?d��0�n�+��������h~��dw�L�\j���2��6k�����J^Ȣ�g���Am����9���ȁ0C ��5�AYmA��Ω��ʎ����6�\3�� ��b���%�.���\�mG�R��)ύ ����S���j��zY�����jY�:����Wh�K�j��H�fw�í�>�3��.�¢�ĩ ��lJ�F��P(�h�cP��`R���"��(Ivh]�N�vs�D�9�6�8׽�t��e��(1�M��
-`2��*�kNSh;���(�#E��nm��`1�p�ЏͫW(�`Hv�6��:? �HT[� ��e��b��)��i[���4q��-6B��)�˖�j�+PZ^�����2C�-���̘���=�>���Ft�����k�6�`d��sb׬�Aa/�Z�2�K����oKO�\�al��f���	���2�9�8�bЄ��v�1����I�� �W^ߥL2~Mۋ��}�GgI���bI♖��-3�n����n�gffd�[[r�gH-�>.o��uR㻙Xm̆n�籓+��V�:�I\��^�Իo-S����>I}�� �N�z�|����?�QZ���ME�]Z�o>�8�T�AF8R�d_ɜ]X����Ĕ�(~#B�P�5�l�`���\B$�sx��M@���_�ְ�w�S��Yg0U!����*������3���w8	��66�a�~�y�"AH���O�kPz��#u�a��3:{��/�=��}���hQ�u�P����yQ� O�;��p�n���n�L�'oi#{�o�ĭ��`�m'���MD�
纟P �{��MKӞA��6܌�0�_�d����4�~'E��j�����?��:�%C͊��ј�1��߶�*:���N��ɀ��nͣm뙨���9�I�	��8��$8��}^��u����@��,F���M��HĬ�`Ez�D�s���W|;E���+3(�bN@ �%N/tB��L�W֍��U��}����ַP�w��0��$�c�GW��n"(��AĬ��㸰>M:��Y"'��>���Fn�"��e��>�X�?�P̓�����J�V�����Y�\A�'�˝���N��/�1
:���\Є�~�����B��sZ퇿��<_�e�i	
�WT�{I�9�>��,�l��p��yB�>6����{)L��T��$�2��q�ֱ�;'�l�;��u3��e��5<�øl?�[_���
��v!�h��ѡ�^RU��a.fT�r��L��w>/�q`��DL8v�Kx��/
���� ��|����r�߄�)΢[��4p�ɥ�{|���%)��?j��~�]��K�^ƕP;�r�5t��3[WT� ���-���b���łd�ρV`k���K�L\ǿ9� Uk�Jɘ�"����w�_�r��Z���_��"���}�����A�w_@A�n�c/^5J��5��(�(����������Cu�w8"wx=�-��ۜ�ؑ��T;B��_8��a��&�Y؈�6c��UGM�/|��M�\��<��a"ɒ TcÝ݆As���l$��]_:���)�R.&$e7�V��O�-I#�������?�9OΫy��BV_g���$O;
�k��|Ujr�)"�OY����T� �3>�v_��Jky�^w�ܯ�d���t244|��Jv(7����X�/n��ao���%�
�/=�U`�&a� ��EN���Z3�L�����V�f�I�RM_�{����ĕ2��\�g{%In<K�[�T����u�w��ԍj�ܫ��f�k�b̯��s�'d�]ɔ~��zb����9� �JI!1�5{d�Ϋ;��L�Xq6779������g<e��8�8�-��|��UX��٬�i7��w��n��j�}|�~�\��MD�n����K2�>�2��^h�/��o���U���:�� �a���ѿM����	�-{���Q�;��Sm��	�,�2570��5�t4�Z����e�$��Y%��(~Ta�U��l�Y�t-�+$���&�8����:h!���^����R��^�֝��ļ����[2�[��z-x�ˎ���3����
��ZΌ.���I�lT(���?�-�a4{� "�_:�C�Hrn����:�����cƎLgv�~�21G��(�"�Mt�ԋ�TI�ʑkK������໎R)Pga�9�?K���n1��Qb�Q����p̯e/W�r�oq�Mrd0b�:P4�6�6Y�y;mdd��u����@�⋮;�M�׋���Y�EI ����wz�� ��̂��b��759���%���+�%0E���y+;�Lb�_�h�:�'n�YԐ3����8��l�ػ��i����,M�Y��ʼu	U�[����޴ �z��˱�qw �O��$˘%1��U�=Z���KyIs\���a�AT���q�K�U����O�����4E�@�GԆ�W7Y�Z�v�~�E��ь(�t ���\-v�h������?��oOX�� 2}d$+��	&^��S�
z���W%��TI6�ݹ�Ʈ��B��]4{��ۚ�������M_�u38��Q����^�X�NJ��_ĝǪrCm�����Xꠧ}'���
�����MnN����5�@�к�S.�1�`H��*B�����q�V��PR�p��NY�"Y�����%���p�"pG�ر�"����,o�$��|vz�?/��b�����S���-Be�4�}��C�l0�^\�O�˝�|(~:�<{�8�w��E�SQWJ��i��e����#�F����e�vg8S{H�L���垹�y�o[��גn���>X��_e�m�ǉ�E��+�e8�,�w�e���D����9�N�%���M�
�Xg��tG\&�����:���S���ZwJ��`V5������`���(O	|�SV>�n�Fuj����l�t+���gt���;#O���6���I)�Q��*=L��7Yt�L���������E���y%��?�;o�9!�N����ּMvL^�S����pӪ��7&XMD�G�0��#����7�J$����}5�^O+�V��R&�b���m,��\+�����(gV�<ɗ�q�O�h~[�?2���z�/t1�)��AeX�U=��q"7v�b�L��ܱk����}6ӷ�Ӧ�dP�s�C���J�%�xv�_��i_R��Պ�x� 4��������9O�rz�?YLa��F������힧[1=(wӇ̹�[��q�Xn�_���)���gq�E��,<�����zP[x�_���(~��#u�����K���?,��������o���鵓��rp;���di�6�uߖ�,��i��'z�_G!J�&Z�&� yO�c �-��C����O�����z���@�jd`0��f�'���&ЕK��L� �M!-�
Ǻ8x��б�lW�ۦ|���$}����`8>�Vv[/������o�a�)�j��ʐk�p��ݷ���UYYu٬�mi�s�!�i
I����NŒ3m�fn8����Lj�r���?�0��=�����0G�����v`&΅�.�~���g�"�n��M�`����WY�.\�I�ę�p�� e��v���վ�/iLQ_M����d�������b��%��U��oD���(�e�1�����oL���9��f�\�FV�`�pJa8�[�R��-��������!|"K]��*''��݈�R�a��STQiN|������p.���]q5�|�¶bv�Gn}�t��������z�f^����ǰ3�.K�H�g-���M
�'*e�*I�̃�����X����Ј*�(1�7~̲�*�0��;}H4fe�z��+۞`u�������z��2�d�b���}��b�;�Y�Ԑ��������vr6��%Ec�j�ülb�vGC����Ǫ�~G����ᇫ��m�i4�H�����&D�)w���e
�!"�H�Kϲ��%p�8��A��Wv�C	GC�w;�b��r'�h���h;�DزÎb)��Oϼ���:��K��<�������;m:�,A_�I�9���J"���}!�I�i��\c�a��G�eM`׹\��F�J<�4�c�O<����`B)g���.m�T)��� U��L����R(����a=���H��"��`�}`t�`a`�)<�F�}A��b��Q�dU�̳v�e��;urXڢ��9�ja�[���i냀�f�ՊLK �T�.EH��0�_��mg��M��Os����G`[�щ�%���@�A2�y�����M	zD�Ik?3$��vK�X�+ևx�J�o�,4�M�Al�y˙>�᧛M�t��T<E�C��tV�yl�gx�/4��(�� Dc�`"o������x�]�$n��Y�'\��ci�w).�,Q������m�4����H���UZ�1�gZS�'�L\�w��H:</���� �=�_h�R��ZJ�$���e�tM�y�b���{�"���k�M�@�_�t��,�S��oרC0��J;��H*��6���A�UW�<>��Xl��U��t�_ʐ������/�&��U��x4�Jo���L�OҀLl�E8u�	]y��v��"����O��Ih!h���R������!=ɫ���.T�����=K�
����E�!p�>��aY
��V͡����1�P����4?��� i�UB�lZ��8l<Y��Qt?!�^�<1���	}/b��r���M2�m*�k���F�X����-0j+d1"�ܴ���F"�k�;,�b��'�dZ��f�V��0T�Q�MD��JA#�#�&������m�wg�ղ7�8G�z������n��� &-Pd�^$+�c���q�W����1z���ҭ�Q/��.�?�`� B�G-��:���D7�*Y���1��RJ��V����ooS���?��$���o@�F���;����˽����������"�G6�w�p��Vվ�Z���HT��¯Y��iY0�%PBŁ��J��E�Fh�Y�T��D�����9��ߺ�n�z-�J��P��`�5��*I�i�<����A ���������eN=�%I��'��n�vi��Oլ�7�/M"l,��˶�5U��cʌi �ϗ�������K��ԇnQ�oB�LD�Cc(�%���i�'��L�A
���a=A�^A�z%W	�{\b����-��)�F��튫�y�y�ؤ�3�W
_�ϐ�˧e��3����K~}{�̗��F�6�Dr)z]�ێ���>�@`�V����I��E�
����[�/��Q��Nhq>s���c@L���[��e�WM��&�K5�,��5�8:f����L�Ze��D1H�Đ�VS��.oYh���m7a"츭;����-��2ޓ�Q ���hׯEgT�O4=�){C<���a	8/�$XTm������R��{��oU*=�w�~��-|��E�p/�1�%dE�~j�}�"X����@L���Z֒��$�)�����w�hT^��.a��:޾+�|3�\}E��J{zߕbnYe�����%����u�d�zY���n7>�a��M��u9،bs��������qe_�ؗ�6ܝ{�bc�X��y���,Q��5����~�*{j��+.�y:P�R�~�����4%�Xc*c���[�?�Fݛd��g�!]"���*
�y^�yDab��?&2ꆁ@ ~���6Y��%SŔ���Zj�j먗:��^k�LX���ΌFd&��(���"ȑ�&4�N�V//wn�X�6��"����p�2җ泽t2�F��D�-�N�R`y�h��C���&��B��J��\�p�a
Г�qJ']"�@Q?#Fܞ�y!ń9�#�ȣ�ܯr�g�`"���2b�6e�N�}eK��sU��*�HC�{\[`JN~�S�[����wR�2�e�I7�&���N�ֻr4�9�|~5��pꕼ���Ld��e����e=�X>ۤ�e�D�~�ڒש�3�>u�Y�iA�x���Ț��Pņ!�f������>��+�-�<-���~�C!�3ud�zLM-E�&��&m,a&�?~���ǭ2�K���sjx�P�Ƭ4�7l_�5#ܽ��}����`�xI@�7$1N=21w'���ik8�a?:��o��)t-s�M��D�F�x��Y�9U�ґ�c�G��*�]n���f����N=܀=�ݡׯut;B��*�:|4a�r�Jv���m�z��d���}M�)A|V��%�ޏ�.dD��(�$G{��C�0�����@c�ckfCm���j�,�q�ؕ��ODW������{�xyʱ��r�t�mVC�Y[[�>�["�����e�rDI�Lx>h�f)b$�
�䄸��P�P	H�Д춵-��JC�@���H��~C�Q�K�2��Y�N�� $�����t$NC�b��i������\����s���N����!4��\����]��K�b��C���;jK�9��e�0aYz٫�/b\
2�D����ܦ�V�	T5J{�d�����"�L{J� E��&�(��m
�I��H��ؑ��_K��5_,s7/���M�*i���-M��n��p�(�F��0f�sM��^���W`	���ܵ(��!f���\̜y}��Y���������.�M���H�y��Z��r���P�3^������×�c���|�U!$��DԄ�]C�����k�Q�T ![��܃H06����5m�v�?��?��4:��{ro''CĨ���_
� !�@�!h���D�*�b=��}���:���v�?��Aod����1�*���p�t�W��6��W�B}���]�Ug�#�@�X$�n{�B����'�����k��Q��L>hkJ��Ǜ]��eљ�.���?�ޗ�ds�:���,�V��|�cǻ@�0ٖjT��&�L��ɆQ5[������ F	8�:޲��~�"Ĳ�HEnFu7��%&�I� L�@�(M:��S����W#��A�h�W�b���M�$D��sM�["[i6f{�I�ZkLo���H}��`^�Ĳ<�#�M�h�b:Ҷ�WH+c湕@�L�Dn�K�m�٥�����|(����	=A�Ġؿ��_�k���DX��`�p��9��[S1�7�Ǳ�:֛�^�.�|Tu��센v	d���~��� �|�+�_|h0ڹM\t�!��Fex"����5HO�(�~;1`��M¢�A8��L\�y�����>)���yg�3Te�Cu���nЅ����ں{n���#�Թ��q��Î��h�=�>Ky�X&�h�W����cIb�ƻ�J� ��"���`8��m�(i.0A(�@j��������vͺ/�+8�0�$���a�M���3Qڪ��a��t�/1�i];W�iVy�jS�&����E1��*�NU�2����.�����|�E��,%$�6����X�^�G@L��sU����ep>�T��+ڊ��/�O����!f�J�Q�g��c�W�UVp��s�N�ׁ�|�(}��`q�����C,^�د�<ܫy��?�t}��7W㟲~^֢���{������>�8����DLR�*�ΟTs|���,{�w�Ͷ�TZ��]��@���q���F�!��h��^/��߽��k�c�$����[GfNS%��,��_���b�Zj�т�4�$�Q�����j��>��?��}͈�lDk��)����|~���0�uob:���.�������[���K��� l:���v=��mۃlN��2Z�k�>����d�v:��c��GU�t��j��]c��	�-7B�M7����?C���pl"�yK��QkM��jO�F�G� �'1b�=�I�8A(a	��O��to����yxZ��5n�o�h�����d��)P��+���|mu?<�Q]XJ��#��b��$�V!U%1k��	�ݻ��lL�`�3?�,ME=>>B����;�#��.����U?qG���c��/��������������Z.kr�*!��$WE�X�[��ۉ���qm�oa��n��[���']�I�AYϻTй��WR_�*	Whuw[�#`;�`:��Ѹ�'p��Lu�9����;&�
�x���F݈�����J����$9��]�$����Z�A^n�il�0~��0s�G5�i�ʻ�y�ϯw�k8�F &��[��n<��M9�s���cQ��(\��0-ڣ.o�9q��(7mh��,0,�!�KաM%�0�-���$���j�Xv�܋S֪��w�z]VQw�9�ʧ�U�p��O�U<]٘WR�w�4ef�'���4Zpo���J�?,c�]�gX��{��>��}#��T��7���
�LV B��%0V��?�j3!>�D���a�k_c�eHs?v�g�O�&��7�$z)�B;��T�������~����I��k��J�Iݎn ��xa���c`F������m+�A��|%\v�d��5F+R���w<���t�"���\�{>@]Җ�!p�\ť�
#oC@��f���3p��B��L�L��d��i'�l�J����ٝ�d�X��G��H��$PMr�69��,1`���Q  ��������oO��9�p��8z$�^l�:�}*K*��{�߷��?��6��ǿ2��:�~56�D�8t��[�N�b���a�2�9@��
��H�@4V�T���7����^�W$�̢t�&�����_�
1\���1��3�xt�Q?�D�W���r���p&(FO..&��9�z)�!>��0F�}uɺ?�?�o*E_�{���1;ܫq��cG,��,���R��`�XII9���a[���-泤eL�K$)$Yl�v�&�PR���*7G��W��F%`{��whr6T��q�0��T������e�+/�~M�D�Ғ�ko�eTb(�RM�ț䟿N��F�]2WK�d��]��3`l_{E�r	y�C�;L�p�����m��FT� -!�7�"�n�_��ַ�h�E^ΨX/|������2��������Q"豞��%:
�)��S�Q9����<�~�*Z���M�	6�=��_B�����͝�ۉ�4�/�Ҭ3WR������7�@��VE��?@��ܖKq��5Y�t�:�<	��h�F�0���&��?��XG���GT~��w���Y����w�?�~z��l�_M����ۏ{�O��^lbVBt_�;a����/�B]~�HG�>�	w7`"���ϭ:��[���j׭�+���׫���紋����3�4�������<���*�,`��_j�z�6m�u�,�q����
x���P�+m��r���<���*M`:���f��D���e!]/>h\���I��/vO��Y�������BvK)؎��Y�΂�C��M�]jgf^����W+:fM.Ic����p�a�_�[��8�}��  ��j#����7� I�[�*I����L"⣣#�#fU&��^dMB���L�*>�L��L��ZX)��N��|hjĎ����E�4?�C��.TO���ȘCm�-F�0Ϋ�)��]�C�6y<g>ĠPϷ�{l�MW��㠶2��w�$�Ƥ_�+�88��V4�V#Z�2��TʢT��U꒤6��a��7�8�� ���ˉ_5�$�!:=Zv�_w�T]KΉ���_	Ձ�hj�k	X��K.z�T<���;Ey��Ϭ�귍/o�ȡV��0���^���\V�f�krg�b��t���aR�����D��ڡf�.z����@���j*d�Y�h�@1QnBvs���HO�����s�+F~�Јj`����8�L?����@Щ +����#��+�dP�x���i��B[��IB��8�{���纞"�/G�ɵo��K>�1�i���P8�N����eͷ|�T���'�Ef�f�֎��|�7A ��7�����t�$���x�"U�:�#�������~��μ����&���}Q��g��;��*���$�VVP�aݝ��xz��<w>��ﶌ��Y���,����b�jCz���+���+B�q�tNU� ��z����]Ǧ�6��`F��d;��������xٗs���}�*i��W󥹸N���Fd2�f�D�F�B(��O{w/���{�!�vb��k �[�zW8�7��?b���u=,?�D=�8�V�K��l�K��}�] 9P�PIZ�8{h�y%F����^�UcZ��E�����瀚���i<�|܋3k�h��C͙>8Ѓ���PZh>�B:iu{�g�% ӈ�#�I�4�_}�����3���8��ҵ��ǫ(��E>a7Kd��N��i>��cX�r���}X�(Os�\��{���lH�zA�	;Z��L�šE_＝�Ma�;����n�ʦvx��o�űD�
w�i�Ǟ`ԁ�vw����}�JЁ�P�ջ�S�$����:��S��̪�����[ ����5���{qkq)�Pܡ�kJpww)Z�%-��ݝ�,����{�o�f�@&���=g�yvՇ��ً�ӡ�A>:.��\i-ч�������6�~�>�|#��B�u�{���e��u��~a[�������X�Kpmwi�P@�<�_=5]����T���%�Z%�h'a��+Sk{,�t�>��z21�q��5]D���B�/&v����g�D�|U7\R,�S������|���';��
�R"�{8 �z��4���z�~j��B�^�-ϊ�f����r�g+� :�NL鱸�G��h�q)ܳ���k,��m�C󂧺������mҏ�P�`Ņ�m @-�q�T;@k��P��B����u�O� ��/�#���%@ɻ:ߖ]+Y�b @��£�
Tc��Ƹ%́�q�r7�h?����e�:�dP�7ֵ�u���{��Ġ����:��OҤO�$}d���-GF��]�u���R@�W�����wZ��PB�3F�m�?$&��^�"=��* ��?��!�ġ� /�,T����:���&���:Ǜ���]� {Lç���@_�a���P[&�쨳IQ!iȸ��?=!��ݪ�eJ�n4����?J 'YY����_<Yxb�bvSu3��MW!�:�]�W��X�[VP�E=\��f\.(n�o�+iMdy��F����X(�a+ÑU_x˔oR�f2�EAj�%�<UH�Ǔ_!o��$;�����Zi~0����'� p��%0�X�'-2jo�_�&M~4�#ʢK�o���L҇#y׻�Kx1u-Ͻ��I��1�^n��mt���6�solQ^!���WS_+n$���T���|%6�)'�f�:b.!�q�2�ٰ/;>;��Z3S�~��3a���M�b�����xLV���#%���ZD\O6mmm�+;=�N͞�*�L�e��K�oc�a�Q&�]���n�����N�L#|����p��beh���)�7I봅��g�;^��QB�K�a=N��}�}c��n����!5[�>YMw$�@T)�~M��Ǔ��t{W%��&5<o\V�;?Op��˱lFC_^V����bk���)�o�Yi��������a�ҭ[���6�y]��VL@d~��4'�h��\���4 ˮ������f��k��*� (rI���ș�H[?4�%�k�.b�q��9@�,�$$Db�Ͷ����S���c���?���x�F�B�4hs��[��b��c��fA<lZe�]D�s� N%*����\��a���3��-2�O&x����F�bj��XbA�{�ի������G�c�}�O��(�J�F*��=�������^�q��毋����:j4�m�߼�/=����w�/1�w�
��7�J�`[��b�8݊���\v<pW1G�\�E��o�`�v�eA_����L[�h�8{�W�p��?�pt���d���@�3�'@a
�5���<��	1d6.F�&ԨMYt|��ס�5y��6��<�Kͣ������+mF��&$֖s�~�?Tl�u�͘ޅ�U��dj�ߨQ��v�T�{վ��;�`J[�;!3"nB@� ����E��f��U��G�AA!�j/�Ȍ�f�5-�g�n�"}Cң��7-�R�/?(��/UfgcUt��,V��}���?h��~y�����&�
�qC�2�4�9�~t&5.߹1�q�%ϨLY]�����$��p!�wc��Ǉ��+���U#pA���Ô{�2g�0(?U=����ވ��4x�[�t��<�s����v�,حLH�s<��vv���;�GM1�晭��	���#�0H_�Lj�ޖ}T��`S[�	�\���~�6���_8������R��	Q��f�Z��Q�/d��1����7�}�-�\/K���$
x�T�=���i��ϧ;�Y�y�e��򰆽f�W
M�q��;�_V?�'���q|S�F=9����X򾇺ެ�Pzi]����:)��~�_3�#�q�fX�5����� �U�k�����*�N͂�d�H�#����H���K��&�I�����+��W9N�W�
��ڻ$m��6
T�����t_�K�V;m˔��3OV�?�#�y��-	җ�c�-q>���8%[�5����հ5�񦕷���Ŧ�@���[�?0�呴T	���)�d[�E����NE��Yz9�_k(���m�^�*�@$�҃����s*K�ʁ��³M+K�Ll�R8�3�W�~��}�X�G��k|C��mAq��5���@)4�[L��U&�z��#F��aJ=ת�L��병O	:�[�8]�m��Ǹ��f;����ϪY�nN����ݵ������-)�H���������-;,2�\�w1�YJGG'7B�,g�[�_�{�D��YT�#���<飂��H�Wu�N������z�`kRO^(�`g�#��6� ��\o�]�ջ-
�k(Ǹ��=�-1H���\G~��*����+C�{�W3m
��#�\N��C��t�[�U�1<)$3�f����\��y%Ve�絫�N�H���OW�J�6��izf�x��V;o�/� ����|nl�7_+^׬��n����)�ՃW��8򥏂�ҍiE0��`#	�غ�^k��a7���	{��=n"�����nK/m0����k�^�!q��[7�)J�& /F����TF�ղ��p#n1_�Ga���h�2̃]�b�\)ac�m�Śh�Z����H�@���G�beת:��Շ�@U�)X�x�YUF*����Eh��B밶=���=�(�N�E�������L-!Td
c�5V͞Yg�3��@�|Ar����o�7����uy�����R(��^$1��K����~����˥�:R��EUv�ǉ!3Z�����9}��7�>�Z�FR��s��s�C)#���~�m闆{]Eq;�A1���z�;n�Q���b2���A�PV+���/�͏N.�Ə�o4�OJ0Q{�W�	��/6��]�5�C�t����,V�2�x88�1B��0}��Y���z���P;������Kp�w�D�_v0g<���})��Gv`�YvXT�HL����u�#��$'"؊K���C������=� s��?�;U��Vّ�|���m�����{y�~<�k�S��b�*��f��-`
Y!\�gq!������F���BTID��Q\3j�;���Ⲫ>���߆0�7X풞[=�7ܴ��!�zRsF����_өw�V|��Y����Zʂ��D��Vg�N�yHM�g�ʡ�#޺czԪ���*tg��'�_)�pQ\C=��K� ;�zъB��j`D��R�^D:E7r�R-q��K�}a��ՋA��q��vV`�<3��ǩ ۷��I��G�����b�����q�17�]��a�p���qlVW��/ED�x�ڴC�p�sn���2���`85��g�p�6ᴏ4; ��[��C.�w�v�
��Y�QtQD�T6���@�2��Cy�@�e��$JGn���)~�ἕ�=���p㸭�Iq����M1��E��CGۄ����M�g���蝡\ ��5"�}i<�R�9��[�nHĂH}���1���{���FiYe��a�M�Nf�CꎓC#&b��z�&ܡ��šZ�'|I��6����L\�Yd>L@|v���x+��xN��Ɩ��}�kOW�h��d�> �׿�ϸ<�4��8�=�'�n�|���	$`/��z*v��m���#��O.��a�E$$R�v(X�#i~tz��Z_�8pF�I�e��D�N�#G��{9�Nת�\s�&߄S�<��r�R�����}�`Z<�nò�2]���#��|>԰;Z�哮�T�R!~ʭ�'��x�Yԧ?2Ɋ��8^o`(�,hz����ƾ��w�NsF���,�7q៖cS�Y{���� :qoٟ�4<���8�D>Б�U�Q�����H��:g^R������"����)�3�r�wԙ�k�/��0�����0̮���g#팱�-�I�#�A��E-�C��xp�F|z�r�IBv�t� n'-���pc��&knYӊ-���)�4)�
7KM ��,nE�]�|���@(2�&��hH��p��x�O,��;�v3�}���|�e�G����Yr��?��n�}�br���C&b����\�����\H�	Uz���ӿa{5X�T�1�玮<��N!��\�ђ���P�;d`��G�J�Kj{�c6N=��C��`�,g�����B����[�B�f]�ն1�̑�z���˶&2��Q��!K�������⛿$�\�0������8��Ń����P{���I<��|R�"��R�� �^�>��
��qgnT��a������[Q���l>�6�� }��u{�.Ζ��m76����kvJ�;(�QWzg8� �""�F=���云���^ZQ~"K�/��	���d@���
�QGX_^e�`#1�BL5��_�ho��M��d6k�z�J�	&��N�o��eƭ���$���i�'�t캊,�D[�� �V�:*�T)J��%�uR����sP��j��-d\���t涞 �2;ӏ�������9�����u�Vv�^� ��}��R��Ŷ�����"�|��g�;V�9�ȧ?�+�N�r(agL�ǘ�A�+cO�\�R�h�����6Em�������c�K ��Γ�7�LKY(E��z�9�%�]~��G��j�w۫X���k嵺xc\\U���ى�����z��P�c��)b2�N�Z�zN�-u2��A�m�|���Mn�݈[��1����r� ������$���MFOꒄI���U��+NS�,0��N�ER�s<��4�5���G�)__�E�	C�>4(��e�!(�_�O�7�DG��$��>���|$4.�q�=�^�w�Wl��j�$���	�9�?xUk)�8�t���0Z��BwN����'�P�GOuc#vvۅB�M2���I���D�1����%qv�-$�&��ӝ�9�?�I�N{n�U��3T���ǈ?�&>^�d�En&�Ϗ�c�Fd	#k���덴Y�w.��A_m5C?�%@8U(ϐ�c%%:���ٰr<���9{�ЪSF���)6���<C�PΫ59�3��w�b�f",8�	�k�ǉ_�
#k�CaӤ�c�&�GP�{C%����������ڔ���쉚�ĦgR
�̽���h����P�7��a�,X��/f��'w(,�Q�_�
B�	����v���MY�j䘙�_�``��N$�Ig�2m�ǖ�@�B�)��|z%K}��70�?���H����9P^��zI��І#����{�#v���vE+���R�8z��sxff,\�dco��z9򧐷k7�&������Z�N�JWK���?�y����4���8�HC琚FԫD|3el����d`Ѫ��1���tw������R�����l��*�s��]L��� �'c�� ��y|M�%��B�Zߢ,w��%'�à\��߶%}�O*7H�J^_~� �@�x�^eɗB�	j ���A������{�{yn��L,N�X����F�{M�%$�k%\��kx��9��<[�>��5�8OW�,��k�cyܥ�տ�*i�����w�۷Ǟ���pO��G��DR6ז�~�����Jl����5t�"h�����=g�1�Ỳ��$�.�����WYMm��]�n{��_�ǅR��?��,Q_GbL��JO����]�+n���V]�L��r_����b�ŕ<f� ,!�dǏ<t'uV���ڡo1�ߕ8��ё���L����Żk'^�*����m�߾*D�c�3�
x1y8L�M��MH �E�=�l)Q�ż�Q��R�b�vL��(Y�d����7�T#֒:�h����9�8�[.*98ir,am
��4U)r�)1`�"HL�u���[k�K���%���w����o������Ff���,���ʻ��{�Pu*�d/��g_�n��@ه[�;��,�gC��K��"��Y�U�vu9F�ʵ�~t�4/��K�B!z�_i5/T�(�������U�G���(<[hÙ|�fw����Fh<ϿGv�]u�����Q3F���cЊ�������P~j4w�:�;`k1� �	��'�WY������(��C��n��f��t+�3����J�0��(,��C�rSe���s��.NV�/�/tU�>�P����禱�~ݱ�"�� Z��s�;�۰�f�|s�]����"�i=�J��5��@+�h���%�Z���ۦ:��}hPА��w��K%rj��,��2�(vjLzό�޶Z�lv_1�}�g���Yf����yߔ�6�Wt���!y��0*p�DV��w<��-�;�C�y��!�=;��4�䭞���&j�g�smޗ�r�zA���ףծ�BV��y��}�+r�l�9�ס����&2	2��*�;J7|ОJ�^�题�)�Ņ�����f�75�D�S��J��#��i\��8<o��0vO�b��D��a95d*Mj���Q8���/	ur2pm���o���;����bZq�K�Oʕ2�v
�;�}z��;y��@D#����z('����s�|��`��IR��z�k�m*��lTb����c^�?���K5�G����Q#��M���k�,�Ctt�0����K_�vTX��y-~�n uT��(Oȓ%Cn���{`�w�|HU�O�>�>�������l�uޑ���R�!ڤ�
�p[�*̋a�y��0���I**q	����ݪ�B��>]��J�Y&�\?̯��8x��ޫ���jH�Jcǳ���S��w���\t�%��Xv���	ؤ�Zk���h�� ��n��B�y-�l��G�R��fUH.�+���J:,�=�2A3��Q�y�Dag��;�a#	f��B�kn9�[L�fܝHڮ��6�Rn\����=����^]N��ON�z�	(���R�֚�x��>���m�� j��р�_:�����|ܹw�zTw��`d��٥�[�[�}p��bo�r�Ţ
A�� �_����+�{%��K�%I�>��z�'��>��H��L��vİ��O܀Y�]�� �]���d�~���A��uEԹI5�8o
ư�d3���@���X7̡F��!�s��3��#��[�h��p@����O$�"�zK�Y$�N&�A�%�[@�Pl*����1j�*V��ݿ�ݘ�b;�����;O�[�]�h�J�k������7�AT�:4b�uX%���<�,:�r����_���u��Ц.���+�ѳ��lq�T/��=����ߌ�꬚y�rȲ^�+�@�kUm;1;�?��4�
�G=�/Ub���i�I\�7��� �mx�
�O>Li}�A7Y�֕���V�z��x��.��$1i@J��#�S#�!�Ϳ�J�=����̹iJ҉e$�SI��_Bޒ����Wc�M��-Y�������?� [N�.Eu��B���}����3�[vl�7�ߞ���q��/��foVJ��q�|Up/�'�& ��nO�����{���2RF������\g���C�uB�����M�3���>3�|/��O�A˃��������B�>!������l��YA/f6�{�3t�k}P�}��x�n�G�/Șo�~�%�@���叇#lw����]��|�'�]�ln����p6�����a�3���,���8-�t������!�"���@TQ����Ԩ���uL���9R\D
�(i�ǣ�ܟj���Co�5ҁ��!,��l��������:���m�$�����v�r�,��������V+�hu����5�a�WY��&=ۖ!\����3��`�f�jX�Ϳ��9��w��H�T0�'9��*u�JX�z�^�����<��eХ�٫�مg�A���&x�4K�A�Ӽ�I��N%ۿ/��ĆS� �i��l�9=��
��gT\$��,m�G>����Li�Ù���՜hL�O���V�E~l�1�}�� _�i�B!�/��M�Ԇ'
�4�3�x]��C�evڲgdY8/MኞNu���f;7��d�k,%Ql��	����ӐA��ܲ�ё��4
����p:jQ���\=߼�c�8�q�Z\��	�;v�f��؀=W*ms�"�Z~�s�Uםro��*���1aeC���X�� ��E���&��sl�o|.�D�ʌi�5���v0�7�ϻ,�����.^�XyG�i�g?Ix�]�5��R�\<�:��ԃ��Z!�
\"|a�6TB��>�u..����|�,bS��A%�Zc>~`�.�j!�p0En��_�j�����,�:�w�w}�M�S}�D"�8�g2�	f��0Mz�T�s����b ��䫅��'f�?��
ِ�O�S3�Gm7��W��ߩ�� �G�O���dn�2�́ATF�W��ZחwH6y@���L�FUp�$�?K�~W6p ����P\SM����v�՜x[:��L-��8�2PW[���D˼(3���S�:� �3�R�y�l�9����1�����l����Jw}�ne�mS��	b��0Ŝ��܀D�.��T��w��c�,R#ng�VI37=��Dzi�gtʦ�`��$(���D���Q����A��68��i��-���9*ĵ_�ݩ�	~.�D���<`��A<�Z�[ً����S�{g�&~�c�Me��w��Fv>� a��7�4@lIi\\ ���X�SV��Ͷ�zN٣���,�̄6@��=e<ZVW�YF:%�AT��9�i�(�g�z$Fa�*M�qP{�\�@�$�j#��ô�oN>��IO��sk~,T샴?P���Z��k`<S��Yo�G����b�S�Yئ6MZ+�0=7���J�GYĹ���]g�y�
X��Vվ�]�4��j����m�t3����01(��|�~��d> ş�0�dp�;�OU��17�ă_��`���(��~���kμ��Ac)E�y�x�.}G?s�:-SEQ�`�_������Vө��Z���te������̝=�͋���8�����]����W�u{�ƻV����G����%f����2l��}�#ΣVbv9�󵈋;.�l9���E������%9NگC,:T���7�d^�w���k�*ͺ�#�5�����>�oLd��c4�'�՟J��D��|�$��4����̌V���+�F�B�4��q{�o���g���5悃ˋǩA�	�Dq���aF����b-c�b��/ʿ�p��g<J�\őe�9�C,���Kf#�������׎��d�h���E���suIh�X��|�pUlqqr�@�Y�A5��ʡ���T��I��{b��lC�S��m���g���.�c
�J�\�85�f�����q�h�iz
����]���L�W��/ҽ�ĘUsjN3�	 �E�j��v��ǲ�ҩ�-z����|�11n1�g?22���T�?j0�&!���L�fF
��8:���F$Y��������t�����੠���C�ړ1J�?���7=���Ό�L���9�$�"J�}ת��QD���ʻ8X��+���n�TW�r���0����:Cݺ�������P6F�hr�DU}Ԏ��b��k�Y�Z�*۟�r/A����}�	��[���c-���
7p �%+�aE:Ψi�_�s�I�r-��
h|�=�B�r,WƏ]d:5�8�����w׾�y����7r�����:�\�-�0�)��$��K����j�����<�)�t��<����<��y�M��Z� ���$���?I:bĚ~����^����.[��'�sq��=#�o�r�V|UV�ڤl-k���G�V�_�f�D�q���j�+W�蠮z��l=!&��L��@�?Q?��C�9K�����s��L����Y����<�Ǩ�wF���\y�f�(M媂՚K�B��3@�(=K�Ҝ���S��w�R"���uY���Aa��8�8�����*�a�d@+q����%lR>�	��������� l@���3!�B.�]6�Ԯ��eI3R�p���ޒޭ���  �9�x\N�H��x=�)�Hn��o����lc��u45C,���&��~��cqXw�z�zQ7h%�
��w�@C�Xo����7�~�C)y���Zq�]0�k�	l���������zN���Z�''��4r�$�\V�C�6���'����t��N'?���Y�+���C�ٌy'@�(�`�]����n�����$+T�`/PG���c��u9ca�^[CCc�0^�σ��韽X#�>c$c�Ȑ.�r�{u��c���b���|�ujTqMmMnELe:�@��p����i(Ԑ�9-�t��>YG�IJ*y�� ����K��"�6�(���!�IJn$�o����|�e��o]��ܟU>Hh����#�o9����g����un�vs�	i���C�i]���d��]�r�,v��~`f������u����G��|���
?'��k�=��������)�bHTI�. _OC�6E����Z뫵���4���}�,P=b�e�=:b��y* ��8�n�Щ3���s����x����yl��4������7_I 	[�2�����:mv����o|rm�����w�
�������Lv�c����	J�o��w.�)�w�=�5���Kk� )B�}�g������3Dw����
_��D5�q�)X q��H�َ؎z�2a�Ҍ����?�'��Scm��
�i��`�V)���}�lfOc�&$�5��a?e�h��!L+��MĿ7J���׻��ݐ�G�L=��2b��_���8��(9e ��b���f��ׂC[��0�r������v�M�X?�t2$_�y�"� You����s�\4��\���榿��8�fe���"�(�W��<=������ml�io�zI�9E4�"�|�	{��M��Az��1}�1��5��mơl�jv>�}�K��#�q�N���])�6�����D�� ?�����������=���EG����]�VX�p���*#ti�C����ON�N�}�٪���t�؜�`m���:٤���1�N�LT��a݇�e��s�IO�>���aQ��pC�-�w݌��-VS[����~+x[R� P���lix�&ix֦ř�B%5�l������e��cG~����z	����w�+���R�?� &��@s;X�w�1���c�
:7k��t/Me��Y����{�t�RQ���4np#6��ȳj��QU��xޢʆ�[�oa�qE{���_�M�O�P.�u3i����'���}b{G����b��n���Q|91�^W���I�I�����ާ}Dë8�'Q�J���Rd%!!�$�t���+"�ݎ�&��f#c������LV�*C��9�X�O�9���3�!�w����l7�bGW��:�R���y`�)����Q�]��$?���5>
r�����M��TN/8��+�����N��-���l��a��X1p�e�^G2E�5���t��ިT翇�-dh�v�K]���A���{�iǚћ��ޜ�0��c���ۭ���^�~��9���W&sC�ӎ�X��j pl�k��� 4��AO/�i�&�y&@S���	��� �	8be-��w�'Lԃ���M�~���H߲W4r�l̍������:����{ai,݋-�m{#-D��V	=�2	�Bv���M�_����M[	sCA�T�D��a>��A��}}�yI>����γ�%���S҂�i��	�z	�X���ςM)N���G��>�g�=ۜ���^E�h�oj.8����>�2˒������E>.P�|Ssh']�}����1�u"8r�����ʬ4M�4痃lam�tV�;�[�9���6橡����<�9�0��{�lfe��;����<ԥ\�&a�/����8��Ⱦqg�'\1Ps��`��)Fl�0-��&��;�$АE;B��΅$B�TY���#L�hiM1v,w�v][�{ ���6�Ö�B6����BV�PʅK�ۼ��W�sBH�'|ָQ�u]?��e���P��o���MZM�c�Ӥ��W;��E�xg�WI����r������Ɋ��Q�Y���))N��M���	"YB4�hi=a���JJ����O*��~���t����z�)d;��X�s ap_�U�UwG9+8����2߰c4�opru��D5���E���"���	`��ky�"��<ݴ�&����+:����\��ؐ��g��)�X949�����ڼ�IF�mWw
����N?�4�M��v�b���t�N����_��֭��W(4�z-#@����}���Q�Pt[�%��zڃ�8%ϵ^f�h����&��|:	[v�G�F�}���XG&.lI�0�R\G�f�{�}2�_�߾}�Y�3b<$A�2�p��H8wXi�˄d�9���N�K�~,ϻ$�mw�Q���~h�ӣ���-���N
tƴ�_^��������?���^���U�y�r{2���=�a���r��qO8�|����� ���a����o�!����7�J���{ay�T���Š�||W����F����4r�2�)�{־����"姯��:+���!���~ E��-�-�7Yr�ʧ���F����%9�ϵ��Ɏl%�B�ٷVu�ƽ1]��T�$R�Ĉ��m;|�/o��>�4���T�	z�|��RXX(�#�i�ьF��t���B���"�k���`��۱��u!ҕƳ����FP,��?���ܫu���.���|��+eJӈ��&�A���v���,i>=�e������O���i�Em*�^�hMV!�%�4g>;�!�x�*s$�Fȓ��[ʁ�bq�K�������� �UQ~�a��\L�$����~лSM��)g�R�����y�H�BX
��3|%�!���x\P����(Y*Wr���#8�xУ�#GKvc,KvRH=�J����(���J7
/���v�'����M�p���Dyp�sI����V�gQT��H�¨���ԣ��y�[�/:�h����	o7ܾS
S׋��b-�t{fQJ�"��W]&%v=a�U�2�ý�e�,3)�C�i��A��]�0^6�M���*�]�E��������;ڽ6���]���r6v��{9���Xh@�>�5���Jb̕7 a���J?ͮ,�%ē{���Q%�x�!�x��?G��*����{�Y�^�ՖJ�XpBg��f���pa@�D��9��RB�KE�V/��D�!(tJ��nQ;��
s1 ����-�B��+��#�8�p��6�"F������aQ��7�#{i�R�G<�ixa��{T$Β��J��"��0쳔H���y�y-��E���!	f�?�9ԓ9�����3}���󯔍�G��P(����q,}�p�
I���9�n#�N�]TdO��_�z�v->z+�k̔�ofTl�da(�UƉ���Hwc6$T��g�R���t����T�����ow����ߦ�*,���\����{��!��r��p�^�,.
����R�bk��� @�WL���:��Ǹz�鐷�Q�:�����7&91~9l��v���Umm���M�~(�� I�V�-�#V��B��䥖<�'n� ����NA����m~�J�0B���p���`}zRUmq�M�s2~a��8rUT�r�/�c�T"���k�<�l�R�]���y=��23k�aYGo:ƾ�TT�s��Ė�Q�/H����iV3U�ᘘ�f���1nbbAo�A�� Gz������W[������#1�V�� �gٔu�e����I=����2fm��8
a5�4d�����6 mR)��_[�:4��<�qI:�o���Jlb��uk�k[��0�J��4%�����?@nM;u��x�%砩�M�p�.bu�q-GS�r��������D�g��i���f��^z5������3��O��\��yb���w_�;�Aٷ���ӓи��`T��A��}���G�$�&���u;ݿ:1Z��2�`�?$+��C�f�_�H��4�'�)��"2�b� 3��`:y��R���;p�Se��q~L��%qۆ���w�&L5�1'J��n�u?z��]RTV���7K��]z�Fg�IoyQM��'*���?����Rȏs��n��U:�>�x���*Y��ъr.��2��g/�Ύ"�Hl��e�Zp{��@!_��sP['kI���q"~�c�꽥;fLV���4Q	�S�.E�wq_՗��߀�R��qY���8z{p����kc�#��ԋ8�lF�d��Ǫ}�FW7�O��m����-$����7��U���I9(@=K�����܀�&�0n�����s��t޹'J�A`U���l$[��<^:��)2Ǐ���~�A,A遁��I��p⩈"��4[��F���g3M]>���H����sf��6.�%z0�`���y�'��"E�B|��� �����@���{�/�@59!u��_��)�C�y.y���zY�xO|e�����P��+��	E������Q��C���%ũGtU, 0w[^^^dd�?��Ӷ/�)�l/#L�".)iF��@�vۗ}Ƈ-M"U��p6��x�g�;���̻ھW���o�^�� ���e�T�8V���I<����vjy��,��~�e��ߤ�	��a	��6c�u~r�v��>��j���$Sm[��D�<�h:�hnwf�l����+u���k3q����a۝�r�E�8�� " ���+z#��y��}t��drP`���^ ��|���p�ij���a(����~
�s�f]$Zf»��R�a?Gbe�m������d9�mb�7:�`	1{�
���ge?�q��T�en�;6"����H��A�ڹ�E�a��O��6�6%-�Z�q���m�ʼ�����5h�8
�C!���6}�~~/�_�=^	�πږGo���cWBs��g�}x㚥bGw�p�{�kG�ϰ{����#%��&xiCG�QZR�o<�4p�z�߷�fPDs4}����\��p�}V���!�2��q&!������c�51a�{�^<��\P~)�;Z�\��T�;�7"��J$�����A'�uԚ���w��+������ ��T���Z�o��6k���V�m��a�.���Oe��*Gv(��m�;�NZ B{f�IL�M5
�K+���_CP��GYM/���Y���5�A�p��9�2���,C˕];H����sa��V;+��č5y�T�R2D<��9����Rֈ۳G{l�in�?��YYY`�J�(P�S<¾��������PFgE������p紉3���;gu%o�F��B� ѡ3�<�ٴ�f��iPم��]�#]���뱈.N��7L��uR�����?QH�͑g��faW0>��$M5N�����P��AQ�`��+��ΰ���s� ��]�}
������>�fFs+̮3��]�p&navz����|r��h��.��\����

�i��BLNګ�z�Zgf	ܰ��è�mѬ��6��&���rs{J�h�kT�9`��<3F��Y3��2����!��V`�;�T����2x��L��Q���f���ڴ�чn�!RN��w(K���`ܞ�%.�,�e���]�Ȥ֟i關q�_6��@��_���X�2���N��;�+f�S~Ȳ�E����g��؜<��sǐ�8�� �Q���i�Ii��	���)�U�4��(����-Va�7�yG���W����ĎS���<��Z�����j.��m<ߥX��O���d���.z0���չ��[���^~6��z	���Gm�s���V����6
.���Vd�@y�,\���g� 2�t�$�12��J��o�O_�7�4��\η�f!�6!�����c�6�u��^�Lgy�I3+(�	��P����-�Q��L
>�96�1K뼱AöEw2��L�\���t��A`��8�T0��PK�I������:�_bđ>�`�O�Wq�=Bhi�C����;i֨�"Lp�@Fn�q�P:��Z�����Uܬv���bw1�<��[�4��pFRLp�qd�G�y��ж�*��zH�ٺIn̚y3Q���i�֛�<ՏZ����p瀕�|j�B���1�z���8.��:n�Ȣ]߂yUX��ñ������l�u�[��61�j)����;�ST=����	;���w##sϬ,n.�/!���D3S�Ӎ�v��������$�4	�
��+bNG��D����+Z��a&�#�?2�.j�9��
5K���fA)�m��մ��b����O^�a�̈Ƨ�)����Ւ���أ\�͊�ݠ���L�}V/����R�����46�]i����%�;z ��(o��a�&\�И���hљPJ&�w^*<ĸ}�BRKKK!�����$���֗^7XY�rN���wY����Bحu�7 �!�w٠�t�K��.-Q���H3B�N�Qc�[��AD�0|�� ��F"�z-��£YL�5eE�É:�y8!|}iڻ����L�s�z�c�:Z���eAg擟v�޷u�����O_�v�}M)������w(P�X� ����
�X!�J��Z,�]��~���f��2�d��=��wם���`snڹ	�;�t�M���|G�pN�T<��U&QLY�Qn�2�9[�_v ���upበtC.���*��u����Ȗ̯X�B6��������V��\<v(�?|0�ܖ�r?emr�:����1��AR��8��ܩ���OVPo�Qg��~29��2�\!�l��	Pe�"�hn��у�ќ{q��稡;i�,�[�Y������+�� ���O����6z����Ӷ6�{�nٿ��K�gu�ӂ�?Q'~�N��3�"3�m'���o�t��(�b�!������ܑh�����^��5�6"���E-u�E�,c����+���P��3�f�����m��W+�$���M9�ݭ2.��T 5��>-V���|;=P/�l���(TG�Q3
�nl���E�6�Im�&H�!~��{�Dl���&~����(Gh�5���i�i��Lz�����%)W��q�k�C{��1mITkwjz���Ժ���̧�D�m�FmT���!g�6sMC!�DD��>�-��Ww8!�leVG�fLX�o��D%���+�C�o��p�LBJj|�ZX�AY����us���o�����צ�Ǯ`����_}E�����CGr촹.ς	���<��i
�kU1���x���1�����95y��@��7UF���N7g3 *w���C-crlX�گ�2��n������j�+Wz������qf����8����a���$$s�I;0��;ȶ�Cm	�+>��[�{���`o`�C�J��G�=?�+fd�[�T/Х��sݘ��ZʣV�f�5�*`&������ԴC6���p�A��2�hE�)l��@���3ؘ�ׄ�Y�~�_�_����U����M�Zsek���&w���:�/��N���x�bf>�Oʹ��^�+���?d�]p��=γ���)��-�ǫY��=�5��gf�Xҗ��Jzo���b�t�~=����I��]_%��!d�� �{�i.dF�%��E:w��;=I	�8�ngh���_��D��:#�k���@n�ū��;W�Z��΋)��3�Zm��[.�3^p��۾י|��~�ɣ�hQ��u��8�h��><��&�r:��{ؘ����JL��_�R�9�蟇��Os�"ȈOk#"Z�"�����	Z�H��]�N��#ve�Է���j1�-�.��6V����>(g�.��#�׀�$�Yi\j.��:	��Ϲ�[y�Q4�[���*9�{�(�Z�B3S&���H��b`B]U H��t�mL���B��Xt�T��'��UҒ7\0�5Gzb_	�dud���ך#��6i��	jQ��=�?��������R זOOG�������������l�����c�@���v�+��U���,�m:i�y���q)�#A���1��hɞ�w�Z�z���f��~u	D�m=���N'h��-ى��a����h�����=�P/Y�z�-+�T;Wv��)�g��,��]��
�#S���6h:B��zKwK�9��YGc��|�;��:&���9������!M��{́޽ő��c{${r�3ߧY$ۓ��sV[P�K��Sݖf�W=��Ô���6{V���m���O�*U��Z[r���e��%�Lzyd���r"W���.$8F��q�ٟ����K�wY�ҙ.O���x ��)��V[�/�>��wF�S�?ASV�*<�,�6���ӝ�^�9�;M�Kľvf����H������Iݹj�o��[�~�5l���u������u��mݛb���_���kFIU<�r1b�a�<`��4�����|��j�<U�VB�J8Ҽ�3�dH�U��h1�4F�zӥ���0��B I��!�h��@��6�H5Ԙ����->�*���,]����h_�u:�bu��f��}Tx�oJZ�&J'�{���ӱ��������2y���?�N���ԋV׭���#�Fj�@U���]�+a��\V���0��IɌ��$�ѳ>��@��
Nz�Nׄ��MY]�3%�ߴ�i·hA�fFFK�,�Dd���K7do1��?B�@�Ԏ��}Tx�<����`����f˟�dq!!���!7���\�X��q����3-��m��hA�Z~B�IaR�fR"ҋ2/��T?��)+�b�|����k�>��T;r���lv�B��/���`�����gk��
>��lg<e�Cr��D�V��5��E=��H;��Æ�ME,�%Ӯ�K�@�rmC,S��M��T��U���L���S�N'��㭗��&H?ܸbF�.עqz����nd�t����X�]˭.v���H ��
`1[��t-X��,p�R����K��mc�����h�(�����qZ�������_�0�@����t���rt>�LNL�f���Y����"�i�=��8怴��
�������A�Ԏ|�m�˦}���_� �X�Z���Pf����֦zi�qL=��6�<Bf�	#H��߸?(�����3VC#��~����W�S�4c�_���r��"l7c� w� �)���B��6]��B�O4bzi �4�^V��;90�~^nkb���2R�~%��b��r)��I	ڌ�os�J���M���G��d�/�T��RR�b$���
���e'�爼~��(��)&@��H��"�R�t3E.(��$�-^�&�f�����b׸��9��S�����OE�;�7��������dP��G^Wb��;>>lP]�U'	A�q����߰*�3,o7�C�ۗ��26�$�%��k�9I���?�a�2v�)}������}�������땀N���bG�}�
���`�A9���.D0)[� ���~)�X�/�&Y�s ?�~��+�X����$�)";*�#���lW��7�`�y�:i��U^I9,�S��<�ɒ�p�/^�Xb��'��ns|]jO�0&�$ ��eۖݻ��4���D:��� ����u�u���B�؏����\��^��%#Sdb��Zo#0�G"��k0>�Ƿ�,w��0���s��c����fסdpc�/"����\9�6_T	E���q��3�gU(k����"ϮV���YJZ���2sT�C�|��[�����x���xց�� A�!�y�����9��LFԚ$Kp6.�ޡ$����*y�)R�znIێ��;��ib��v�~�9^t���{�Os3��D�*�$��)#�T`���sF$.�#Z�zW�H����8	=ذ�)�_ �K�?�n���l���\s��r�.c)H��Rﲧa���^��2ig���'��f�ң����e'�;P�їd����v�_���Wv��+���6
�S��&�Q������?�4:P�ΑIEl�	����>X��վ������=��Y�4A/��63����3�*9��C���\�� D �#8f$����
��޵w��\�ztG�)�e ���f�M�P<]*���:���8���m��̊�o��O����1�K��O�q-��i��#U��S����p!���_�Ut�/����̍�"h��!������}p��}�b�Z��'���d)��@��n<3
�~̟�3�ʲ�j}��Uo:�[6�����l��6�O����vB���H!�w�5��s�΃@���.��!t��ￃ<;0��l՝*Wt�S7u|�1�:l.�́axd#�ɢ�&�c�{��?����7�6`V��㚑�����o��8V��q6�W?`��eWd���P���꛺Q�Oħ�����q�0�� T�k�8��{xMk`�@3H������C��ͷ�}���
��-"����CJX����R��X��n����?��mo�b��8��#k+ip~~����}��K�a�QE�s>!�<A��*�_�F�{S��N�9�x��ÿ��s�4��rp/ԙ	ˎ����Zj+�i�Z�����ڒbJb��\&ݜ���X:��agG�E=ݗ���z��f<��~�I���mc~�"��������ZIh��%�w�zp�_�>t��K�����A��۪��T7���ʹ@�������cF�nݥ��d�^%�I�K�l^�|��D��d�U�BZ��:�|�[w�A���Y"�q�H�5Kr�����t2���c���pQ�2_��n�턘7#ݶruu(��v�ǉ����o_P����%��D���:n�8�p_2(k*��w\�I��_E��A' �矛D�:y����+b9��[�gLFG�U�4S���!�n��M���A�SY�����KǚO?���ki`���s���Xg�@C�������8��Up)E�ӵrhp�J9A�4�����_t��6�M+{'{����o���&Ã����6;�X���5��I
�c����ik/�ȓXdY��I����8���Cz����� ~�Ҽ�Q�N6��j(�D�~ن�4��Ґ7_O�/��{��ap��\-v�=4ۚ4��Z%�}�`Jw�����\�W�s~��S�frٌ=��Zn��q��.���6���b���QRn�?�p��>�0n�����bj�q~�
S��^1���l=��D`s�����&x7�%ν.�
���4y|N~!��4�� ��M��QeoQ�p~�{Alk���	�MX 1��v��`���H>�G������yԅA��zgpu�b!��b��22Ys�.q,LH	��@��QG�0E�Pt^�ӵ�k�=DN�,��T���恑���T�z7�~�}F"EP!.�O2��TƕHW7k����1-�c���~W�A��N]�;w<A3�	$�)�
 H����#�1��������bR���~33�4C7)��}[��_.. ,�D�^@� n������'�<�u�������߮^�$7U�Ys���ϐ��3�[���=�i6=������l�F��)BPWZ���~)�����?l��%�4�|�V�I o�9ߢV���b�
��i��3J5�^���KZy����HV@����-n��3��q�p�±����7g�CW�ޔ5J�Dg?�o�7ۤ�_����.(�����Oګ��K�a@F�+b�tI��L�z�G'��i#4�xkύ�E�R�ã�N5y]VG��J�N��S�_ ���a���7a�*΋3C��,J�ښR,�s�y�]@0��o��_�G��Tp�:���3����׾�&���[�wr�T�: ���-��S��_c�1�ҷ�o�<h����+�9�Q�r�PP�B�9���S&�ﻚ�&cr�-��O@K遬��j9O�=[?�j��	���q���3�eTgk�Ii�kl7��hg�q)~�y4�����i7�HS$4&_�C}�����F�w�*Vș9�e��{Z��V�������^g�%��i�&�Ǣ\��s�E����������%'�gsJ�5�/��z������5&aIQ1���>�5UP_݈Wj���o������r�	��t~������Ҽ���c^��b.�GU)�$�͛Sa�r7(�K�n[���'s�o�_�w�F�L�`������h���V%�!���y��?�I"�\,���{T��Rz9�V��o�-��q��t=��&��jm��k���&�H�<۷Mt�lA�q`����y���p����\�z���3����\������l���w�Ŕ{�RtmBV�ƾ���k�ə���:P�2�A�~J:j}_��d�;��������>�'�A �h�bss�q	�~�2k���2���]��3W[�n��<��z/���0�d1a���|h�]ck�o���y��-�K��`������&�J0�
�5!T#�)��9y��N��ɭC�dHs𻥩'�GL�Jc�����ip��cB�\(��#q#�mi��J!�qԻ�hW������U�0C��o�N�����y�o��O4�},ú>�d�Ȃ���z�yQ��L�<9��oK]>j9o"�rm����EJ�O�ޝ11����oe�����`u�OaBY��us���văl^�1a,
�<h��k���y|yDA~���%�ON��n:�ݵ+��mܨ��|fȃ�K�s���f�֘N�MY��%]$!W�?,BÜ���z+�feMm=��)z���?W�%<X߭�����%���gCC��;�wT�ؾl.0��P��k+<�l�PY����P� ��Z�G�7I�<�[�:�`�t���5c�}�4c?U������2���sD���㕪�[�QC}ݨ�3�G^R{��ͫ���r�֗�X?2���[�#8��M�뉞ku�k�wܑT�Ft�]��vmJ>~�J
v��^�<Y�IԄև�̪�H���ɟ��ƫt<6�����5ײe����3A0PW�F�Ҝ��2�^Dq)Tt����eI�X�(#g@<�m���QR11m[�N>�7�BJ��n�"E��T<m��c���S�Qb9`����O��LM�I��I�A���0�Q�����i�/��k{��2j������6X�Et)�kW|a�Ý�������{�ڔ2B����#���N�8Bv�n (�i�_�����Q2ޟgq��HB����պ��'dD��U���'c䃙�a�=��򺅘sª�2ƌ�M��h��Q�s�Q���-��:#���sE�����q��O%.�Y֧~l��1�0�#=���WD�{�v�::�m�>:*�sIm�&%�!��-�%��YN�!�t�����H�mWTeqr4[�K�Rq���WL�=x�VV�6	t4����n
��[l��Fv8z�Q�?���5�M_�=���%�Wr��҆k����#�l�(�Y	.�ӷ��1`!���b�H/��e�m��/%��֧>���L��E?�W�,ζ��7�BS]�4L8�Xtٚ�,,�T6�q>`�w�n�HB�����ș�/]��[��w=�-�~N��ri�#o��q�]�e���E>��(�<���^��c|��k��w!ۿ��;T��s:i���5i�l�/���ɺ��u,�xu-����<M�2�z�ɏ�%��Y��7�P%�>�ӑ��B[U��9�����`V�3s�$s�o���w#�$䣐�,�׻6��Y'\!� ϊO�-���y>��w�U���G�D��[]�_RK
�)�ӥf�f�FP�,�?���6��x,�܈ <��&4�E�k7��jx�.k�@�&��#����ՙ<&M-��w�cK�>�3Y����`w�6C>}�a����ugv�.`����P��w}�)�˃O�Bv�tͬ��������_�ɺ'����A�:��o�y��NeE���T݀�S5X��ƻ����iƾfu~�@�����<u������2IKK��_���{mB{�6��x���~��k�
�� ��5�.<r;=��&��:Y��9��I�x����CnR+E�m�61���������%��\�v�������U1s� P���8U�[��q������~/�������Njdo�g��8<��SB�r���{��@[���� ����?���j�X�i��z�kt�_������
���teC�#[�7S���1��O�|�S&x1jm�c�yZ������Q��B�3 G�OA;�����X�$�hJ����T� �z�V&��9���Q8&��1�:P�p���Z�<v��t>�7��]ko�'�RjBi�u<�E����l���
٦B�Ts
���^=�=jM��v�����;zbd+�lJ]����s~�I��~.V�k��+�Ԛ�l7�\3����.c�<�9���0x���qŜ�����x:/�r+���%y�.���ￕ&�R�ؒrr��,,�QѨںڒZ|���U���c<�ؚ���З8�^�e�[��p�Ѷ���5fE�e�����卜N!3�t!vQ�`pW �֏����S�,��Ʌ%������h�KK�_h�R1�ejVo�<O���t߹\/yX�M���loE[�s����R:�n2�5����
�Ey*�.3=��y��Yjj��diT�[��"pQ��3���6�z��T^�RG�E&��d��N�V���j�è�Jo���bs� 1�7~��7�ـ�69N2��n}�ʠP�H$/�ī���ɽ�h9<P��n|���ooK�V���	Yuݹ�V�o��LE� e0n�7�18�k�*Gp�t��PA>?\y���m�9�Fl㑗�C)���q��"2t��Xb���i�=|ﶶə�P��#I�I*81������N�����}��F29�t�W �bb6�vr�>o��> /�j����!݇���]�].�HBw?{�.�^����0�?�9������Zym\�ڳ�0A��+�hȠk�����j���M<�[l�i� �G�<ې� ��_	���xT5��H�X������0؅)��}I%�yGKK��T���/�R��,)f��1�e�r|f���L�IC.~I�$k��O�����rG�����$D-���B�h(�Dml������R�=X�eqab=���[z���n���}��pX�+~��x��������j'/D�q��R��7f��M��)���G��f�g�s�ޅ���=۷}��G�	}_~��`��BZ����t��,?v�ɷ1`BR�.Nsg�˘r� )����~����3}��_տ�vj�E��Vw�и�^�z��FI��:�0zO�,�z"u���hn$�ĿQ ��cQ�+a[[������}�[J����H������р�c���{�ِy�3�����L����`٢���I��)�ZѶ-z��o����^����ң��·
��Dc�e�TD��j�Q-��H-�؏��j����Qo@u���'W��D�k��Pj�R԰�������a����(�C��Ad��w���j��xQH�U��RDj��*@�\J�tn�}2fD���WXI���+�>^K8��9Ҙ�5̫bb�@dK�%���A��I{��!�h��8��ډd|�dۉ�%����$H�nԵ6Y���m:k�:r������ى`��s~�Dy�W*2�Y��U?"C�B����+m!Q��nnn���b�w�e��Eߛ��[���ܽ���	D|9=$6���~�������+OG{3a6�9 �ؿ�s���<�:���1yvs۠�䁈a1�4�����a0Tb+�D��	·� ģ���}U�#����éA���r؄�O´Ԥ\]y^:�v��r�py_k3IK&��E���:V"߁f:�%���z�LD�Uj&M���6�>���f�k��nsU�Ƭ��Y�� y�@�#������%֣*��6�vB�����N�֚�+��������9��� �F�-P�� �@O�0��ӓ��Cqa��H�A�ȄM�]�E�RO��[>��k�R���f�Z5<��p��B4T��IH<`Pe��{G �vDX�jwEA~��{�ܑ�J_u�;���0X2�>��X��D(^A^(�ݩ��闫FF���Y�M��x��?�~��	łY�kD"���y钥Jl��\���)B
LG2��)��'0^��j�x�G8P��Ҧ}28v����1�{A����IFJ�T���@BBZ۹�^���4���� ���p"ŵ� -��T����!����~�>|47UI,�m	�C����|���$� G�m���>��;��XF��S*�������&�У��� ������]���!�?����EoVC<w�<Z��5���ns/��г�����*+��{TM���K�+�z&�����'h�l���:����&���_u�1;���2����Q�}2�@C5@瞴���k쨨���),�C��:�~qqaz2��;��� ԙ546Z�}%��m����mhj2�.Q�m��5���@��c�0R�+$�W�� 2ۏ��oн ���`�\��|9�BOW�t�m�ԭ�EG|�jʔ
�X�M+�� ����f���^�ڬ�e��W���L�+��XR��zH�h�=�'5c�{9�����A��[���E{
9�"8�a�/���.�̨�*�؏f���H��,,���=:)�:��KR�̩+��]7�SVs�5ɬ�����W���;�Oe�#M���W�-��k���BLPo9��{Y'Xq��8K�;�-��pZ[O��8�^�����-�|����	ψ���H�~�ֿ�ϙ_���!�r�{�6 eˁ�0`�I�к!������թl�h��������3�5���+�����s�������Q7Sm/U}y��t�Q��UPh��[b}�u�����w[e✝wTj�"��Gߢ--K�9^K�V{O{�C�>/C%���v&A��.�R�$ta�a.��Xr���
j�Z"����(�j�������k���i��֥*Z[[[/G��X��CD	�~u(��s},��*a͚��G$L�7��Ԃ[�l>;g(`��bw����֔����y,r`����1���\����y���<�ix��M����+��nŮ��d����Y��+����ى!�h>�Ǽ.���@�]��g|NN�K��"�UTa�6�AhE��
#�hDe #K��}G�t5d�}���R��[�Q݁����G�1c(a$l�9�ts1/�����l�[��||w^�'����p���p((�]��,x, �99�hk"}�U'@����t��&(�E���ϖ��88��uk2.Կ��:,baa��:���� R]����"�����Q���n:� �t"ZՉt�'C2ЇP��ֶ�8�G!��R��lmp[O��� ������o݃i�A��:{�6��cҤ������P���nӐ|۽��Rot; �*�@I��Ҥ��!ߓ�j4�o5vKQYd�M��,W��ӓD]E�7���}�-�����#b.��g�4�).�M��:�FB�D���±�Q������6��ѳ`q�QPJ'�~~J�{�=��3�b"�=nLs���<8.i)�DO�9� ݎ
er�]>��[�,�B��#��o�[.w��;�����$�ߟ�f��E5�a�G�-�m���)��~����}?�|IWz$j={�_VZ��Z9����N��5o>���@��]&��6q�%$�;��vt�uIc���d��0��cg�x�#�|����mh���z�bd�Uo�F&����,�LČ�P�`k5���SmG���ҟ՝Phjz:��d�/���0����t$�����KY{049��_aޒ�'�'�xOw4��Ki������`����r iU�&�+G1W����U����� �+�e�܋���cQ	��Hb���.wG8�?�­5D.[�b�B���s��Ė�Ի����W�W��@퀖zk��N٠�o_(��g�(��g�{�3��A�6,��8V�8DA�\
��G���]<�]����	�p�\A�f��~������^����;��@��Zw@,Byhd����nt]	�IrugN��tS`C�x��gY��2,cbz�u�����ܳ�yKI�:x8�vg��V���'79�B(6�XI^upu�Ĩ Гk���>X`Bp��C�2�Á���K��5�����D]2�RM��u�J��<�1�f�aw�� �S���kg�'`_�nu&��e)�/�U���GH�iao�!-�&��_��)���h�q#��BgCl�	��
��@r<zy���Ef{L����ME�Ҹq�K�,�䞣w��]F^E�(�U�b�𤋮���Í`��`�����|��������&Я��0c��2��3����}*n���K���[��x��WРұ_4O@#��ӊz��S^�5 P�j��CD3=�;Cz���*�xߪVM4P���np�Bq��O�u��)/�)OT�f|�@�R���-Jv=�v#d�pW�� � %?/�VA�u�.����&�$�`��#D3�P��t��㊄��B�1�����́�K����y����/AaYș8;�<��[C���{|�uύ���x����l��r./��H.2�$M^���}�Ŝj��ٶ}�IYv�E:k7ϳ?⒱�)�id�~�������/���lm��`
z������q�} ��8���u�Y�o,}"4AU��*��Yn��,6��^ɩY"�^D�3�Q7W߄.���9.J��Fs6~��:j����UV���V���[+��ot��m:�W��M��<�E띉�b/�I�S;#�J�� ��\�B�<'�A�ir��Na�����煉l�K���ިפ`Ѓ�U%BvE���`,�8n�W��#
߻�RO��)��H���y���ђ]Z�t����n-��w��)2��W?��A��'����^�Df�����vh���P��K��λf`wЉ0ܵ�
�=Rts��2a�r�g6�ϓ5AB���6��N�	b��B����r�n����/7NMvH�@&}�lL_���(�
�v�-��2���L���]5̿bDV�]�_Q��с^Ŗ%X�	91J,I����Ә��_Ϳ,�X��*�![P鉒�t<���gy���|��Y�s���(a2jh���9( ������M]4A��B��s GuǗe$�~��ٟ����#�.��c�$Q�O��"��:e��ۍ��;�M'���+�+�wگ�yZ���&�|��X8�_䉼~��ް�v��xTn�3�[9hq6�̇��r���� '��X��I�L���W�!�SDJ?ck�	mS��\�r�[�z���(���eu����AFLr���k���[X=�q�0ø�c��H^�v3=^��<hĘ"*A����Y��_4��%y�)���L�*�q�m��}�n�+\�F�����Յ�|Y�k�(��n"�Q�Au'E�)�$ "w[W%�8u�����Xf������LIG�WM�/�#'Q�ۊ��)D�� ��\|�7�T�߬����r���L��>�,y�m�Bs���Z�L>k~l���oL݆�6�@�9�~���Bd�gu�q�l�c:���3�j�m�c�ms�QLKo�����'��&鹫��O��"�u��W7�ޒ
�3!��U����`P����$(�ԉx�򡨵
�mvN��:��͸;��~�~��@��W`���t��W
��.���E� �
&��G�������:���vG��u�U��P!Q�ޤ1M)!(��@���Ӱi�>Z����D|�_�Uݵ1�2���і5�&����]�}�+>�.ح9���:��N+�Ԍ����x����p���ʐE�7������P|�8;�\�=���0����	���Y�������3P��VÞN�k�N��K���F�W!zЈ��:8`U>^����|��9913�e���~t��%���R��J�|�] �u�P��ر{�������� �����C�in}mG��������y���/R�2�_��>},+���Q_�#������N���j���h�[LbI;����݃2�u�4Jo�nsʜϭ���ytk��q��g����7p�xU�,k�%'����R�%(^nJKy�	4�1}Y|HZ)WM����n����@.]Q�"2��Դ����=:�LI
�����^!z�~R�̟"V|���U�.grwv��8,X����?����ִN���[���$ʒ�H�yR׽�`53�����5�p�ӓ|7�s��z�m�����i��p�`�g�U�|Q��0�8�@�c'�F�o5����pWӑ?'��]hO�Tg�����1Ϯ?���0��޴~7�h|q[s����m'�p9�l|������k6fV�3����h�A�T�&)���`�	��f�ۣ��$�IcL����:0ȷ[e�Ź����0A� l٘;W���n� F���]Ȋ+�����<��v��Xw�R�J��SB��	R�s@K�]��'�~�T�H���]�Ϣv�d-C�.��j����j��k���}�_��Ү`G� dac!:��XTB�?�ţ�Uh3��9N�5D��=&��/������-}<�5�Zc<��9�*)a�v�_gQ�쁩�ǁ�#���icJ����$�"o~�����~=��̡����!<`cv`�z��?��"�X_U61^:��w/5�:��y��֊���tл�z��朊#oo�ɖ��86�\��0���V��C�wF޵С�D������yk52���:�����*��1	bB�S"h����zI�P[iO�����E�D���/(a���w��Ƭ�g��tl�Ӎ����Y���ϑzH:W��6T\}	"�Y_PR�����)�g{����AtA���U[W׼?ՖHScW������xU�.�	�<o���
I�ֈ��**��t�~-��8ώ�
���� ��Wf�c��n�4=��"���*XF�u����[�$����~��\j��!j���TLd���(��R2���΂�~��ɉX	�t1[_'�^(�P�M�Dރn�)܁�{�Cz���`�$Cm-��TW\�8�z�16��!�Ђ��Qv앸��"�W��,nn˝�A	��OClՌ6���XȺ�=4�q��x�i��ZΈ���:-���(H|}�*K��l�a؄��1�((�-e�~�7���%�	�:����@�Tc���8h�7���E�lXz�
���r�Y�8f��+1��n�O�$2D��~� �|�/��p��K�CJ21_�1����rs��^q
��Pj;����j`�_��닉�E�G�i%
hd�uƐ�	��H��蹜����-���Ⱦ���Ͻ�jW/�}��oNܙ3�N�7�ĥ�$o�,o>\>E2���[�Aq�0$3��Ǒ��1WZt�I̋�3K��|�>6]>��=���Cw��&^���ZT��?�H��Y"����S����]�7Jns�+��C�-�6A�'��FF��%�f�ݏÐ��P����W;T%���B4�:���Eo�'�_�?�.还��~����r�1(���ɻ?='�����dm�;���U�lY[�����m�?	1��G6~��*z��o�[�}���pq376��1Ŗ�ª����"��!M
X�E~D���Z�e)�y//j��/ו�i�U��ݲ�jH�Ռn����P8��M��ʪ����'�כ1��*1���A��=�4ڦ2���j�F�}02�7_g���u�����ii>(�rO���0�)ҽ����9�&k�fub�ڠ�8H���ᜅ�,���Аt���5����A�JNx4�J����)��r���Y1]���va���Fp��A�<	))ࠪy�A�6JG����w� ����rl�MlUVxx|�)]_p�?�U���!}���W�]~R���@�7a>�T;_zQ�Y�2��.�?�_��������Ø��z�&q/p��M�Z�h���tTP&0`�q�n�9�.|���� �:P�$�N9n:>���`v��0�W��B��Q�[Z�y�
k��y!Wf}u���8�馉s�
� } 1��ݽ=)y�c���"����EL�Z|�,XP.7~�Gy�q�gu9s���u���7#����H�-^�O�������s8�o��$��!f5��qyh,��a���W0�+��M��R���I���K���T��ddrKKb6���CE"i-�]B�0�4�B�/4�{,�E�P(��O�X�Y���Gya�	�U�nK�c��ۇ���,���I��ek��Զ���+�E�'�$$�G�����|��8���7�W���9�,�hi�䷥qh�HnӪWgs�>6,�ik��[d�,�cHNC�rG��z4�DTa���OX�S_(
j+��"=<]UD3K6��{�ַ�?ؘ���Uڃ<$b�2|�-"�6;��,�KW}#��C$�Ϋ[�0F���q��P���-'�{�)�NA�yE&ވ�V�b
��)���6��R�6t�<Utii�����Z�t�!�O��{��ق�����&c"����Z.t_8������aV7�GS�(��,fTo@<�l�Qz���K�����:�f�S�ӛ��jE����հ��1�㎈
�|� {�m2��,Q��4�H�0���xi��+�f��1cϣ,�GU�uڼ��� -�F�;<�I���7���v��Q�/�Tک堫٦î��#�q� CA,1�~�B����%�a�>����؍ ����'yT�[A��"p=���ewW�r+�I�6TR�
)Z'+���b�����K��q�8�
K,8�t�V�A>�wz:J��	�82�r��q��m_#hҙOA�����;��k�d��F�[8���
��޶����>)x� 3�]��ǿ���>�>�S	v������LN�П9�aV�	����:�̃`�%FW����4AGG����aO6��r�	$aџ��}۷h��NR:˵Qk+T������ފ�u����c�T�Z��Qt�0ij�l�w2vv�e�WėY¹�)��H������i� �3s����Hc��f9>�#
���A��/�L2�C���q,L�);�c̉����@GC;�E�����j,�����M7eU������6��}�m>�z�r ٛ��[�E1�a&<�?��:*�����S:��S�.I��隡�SD�AA��ia�!��!���{���5���ଳ�����s,���·�ArA�7A�?ҏ��k��F�X��T����'d�Þ��n����]]</SLL��Ŭ�$��o�&����i���[Wv�"�Q�d=K�
 ���/݂�1�ۼ:|[ǥ��W�v2u����u9Y��u���w=�vࡪ�W?^EU���'Yk-��\]��sw�Z�x�|�@�����;{Z':R��~?$?�JKKN����P�@u�޼+���k7b���#�h���OMV��g���}�viݧQ���@1Gl�0���-��ڮ���L�&;	_��p�nl?Y��-�]��/Fŗ�������s��OKio�U�;��Z}8�k�gn�ך~���DZ�h���j��*EHb

�u4I�c�&��׳�lmK]��gA|�+��BGG�ւ=r�9�GE������3;4E�f�ŕ��ۿ����1�ϑ��$����������_
!��&���Fh�Pq�R)�l0���Z�u�⽞pu��x 	UaN�ñ�WN�$rZN�:V��y �p�!�ig!�0���G��*���Δ�јe�ϞKp�͇/I�d�c;��	bEU��R{�C�kB5�Zx�Z:��ӌ��v�������-��.�V�B����"�u��9>a�zZl��{:�-��F��Ġ==���.������]�YI�?�����Djk�>'�@/��ʂ	v��/�����X��U
���;��I�0Zt6�}��w-�dq0���m���/�ϛ}ha�4sE�Eg���V_.$�4٦��_��*1[�=�o�Q��>���c��P.W����yj�2�NVv���b���Y�W�/"E<���L��&4p�w���|�L�Th=��!��C<�@ ?��4I)�i�r@�Ԋm�}��{��� ��f1 �d�$D�~����H�?&���,�$����Í�d4ùJ� #��-��E�?JNK�Wd�s�G!��ݫY�[ſ�Ԛ�����fP�LS�D|�}M/r*�Z�uw���v��X�ť�njW�Ly�Z̨����¸���紲4�ӑ�"�vg��|��e���L���Svb�߆W���WP��oT+��0rj�*kj��!����[�����A0�i��N�Z����;�^[��Gi�N��&雗�~�T�ߧ$�>\cz~l�lזy5_��w���	w��9��.S�x�$4�~E�Qa
�r>��h�4��܅�K�*^b��d�?8��Tֶ����d>���8�&��3�>��2W��vvj�Xp�!>ٌ-�oO���'���a%���10��AW��$ؓ[ �,����%��J7[t���c�YAi��f
+(�*��xr���6&C'�)nw�}^�������k�$��_2$�=�%U�������1�;�1h��˪G�O!fy�-Tn?�c�&�&��c����6��r��)_�hSK�s����Aw�䃣_�xS���x�˵B��k6�3wyRHn�^��p����^�����u�'��5�K3����+��;k:S�;?nV�X�fB�����S��90�Ԓw�@17�t���^�fg�{D�n40'����WVjv�BFh(:#���$�A�:��ظpwC'2cu��̚沉����&q>�`�JAj¤��F
������ �9�	n�$v��g"m��=+ޏm�+s�������+��OE�W�j��0g�WQz,*��b�ϕN��
�ʰI�
w���G����gffĭ�h��^�9%#��)���J�=�f�N��6C��d���?�����E�;̐+�� ���4�8	��3�C8Ҳ;����F|���3[(ޟ\������g������c��^���.����\�=��[�rov���(�����Au)��6�d�Z��N)� 7MCl��� S0%�Ve,���:�Y��sa��3��L���{&��ߌ��{v 1q��ʼ�fܴ�]A��4>ԉB��r������	�	��Α��>�k�6��f�&���^��:���V�_��Yd���h�v��N�~�6�da+�j��.o�����E��+v���k��Si�8�r�К�P#�������r���+�Y�g_���[���Q;ntJ�g�)?�gǵ�Y�.v��c}�C|��ɕ /Z$�Ci��lz@A!c�����{՞ns�r%T1��״��pW36��<�g\IҼ3u���t̃�t�����L]ڰQ2�ݘe!v�\s`k)���(9l�Z6Y��(?ں����iZ�����Z�7�Gd�}�ж���JM{�y�'�D���"��=�\��f�`[k����{��W�Y�<U�D�~�������z6,����n3��� A�[؅<7�+�ܕ��=[�
��<�ʥ���y�*���i�Eȗ�zng���g�#l�pz�2�1:Q�$aX'Κp�k���=±�΢ҍj���U�P�� +?,w�!�ɋZ_�����N�����	�.���n�W����4�����2���>��\����=Wx��FQѹ��hv� �<�6+I�a'U���,��g�sav"���{F\��b?�*��{����[�GY�e��pw�����1���n��N�տj�-jƂ�:���-1�1E�G	�ÁQ���e����ʆ�w/�-��0�q���V���:wa��g�|����y����-̰r���t���`؅FXy�3�����sЧ��[�;��X��Hk\�c��>�<=ۭ-uA�1�I�J�x5�a!U���՛{^�Y�e�3I=�w*��.��i�?λ�Af/QY�7�%3~���yv5I�[W\G�$s����4�~�RWUH��0�
WCZ����G�������̆[Ƨ���	�[i�-n�GxD�n�*��<u�H�5�\�;�\	�{�z�O-6Em��j8��i��ꍍ��7Ű���͐�����E".�Ń�:TdCqdy�����9�2,����'_uǿ�TT�H.����_�+����}��Ӭ��_B�յ��4"Ʋ���"gB],1���x�'����)� ��u���)͹�Dϓ�5Ӭ\]�KO����%�YM[�3�	��)G��:J���p��L:��%�c���Q5"�9w<�R7A����xn٢����"��+Ո���5f���@�8B(b�2���p����6�o4���\���@̪��/���<����f���w&����a+}�h�ڔ�m_r�I��t�%��3hG�d�Z��u�p�˩�2��#��ۻK K�>�qK;�D��&�i#$�E����V߭�'��*��*�"-���h��t�A$�pC>eU����p��Ap*�{)����2W���*q���3ޟF7[?�O	�C]\j��t=��6����ͫ�����X^k*Ə���,��\'c���B��M|��ZJ���`as���'\�nwvb�F��/<e��A:��cU@�2��=/�g�x��~2��8�ֱ:a}J8��g�$��)�����m��,V
��2}�'���b��@=��om}Z��έF��F156�[-'�������}2h\��?١�O�00���g7���!�5����u��b��)�+�$C��c������ȓ�� �ZD�
�#�g����Fr/��u���(T�:����s�p�[����ëa,����E�q�7�$0j�p��H����
�Ȼ��OZ/�v�*W�^��5�[�B���	�6���"z��cR�1��XB������j��l�<�� k�/l|�t#��W�͎�,nV�y*�
4�Xlۢ�$��U�m��}MC����_\Ot��������>��g�`���b����_ʋ�\�ܸ�ǯ?��Hx�Ny?dڞ��Wu�|�Pc%��F��;f��.E��ty'�Ɔ����|D�M:�㔗�_�e����$�I��+���,���̾s�p���e�k�$:|LT�C�K�)��������o��.�| �flՄ�29o7��Il�����s�Ћ�d���zM��R���?k9�'ö͘�$����M�5i����[�����'�?�@}��m�w���K�lbkŹ�w�l.�'�A�W�?�S���>�?�2���0^<���%E:O�뭁'�Q\%�%��j���x"�R{�a��w)��l�.�3=ny_��H��	\�Sz�����7��Ч˳��\���,��Tm��f,���V��M2g�p2[�'�������
�N���Ob�/��C�/����k�3����>xŖ�3���(����e�����6�3{4J�/��h�iDy_��ʈ���W5��9�X���D��7��2_��h��@;�hh�9�*	`E��@�X�|�H֣��+M���1n0��͹�H�|�E(1���v�����n~��D�m��Ʊ�4�;�y�>Kt1N�n����=+��Ý�e%Ohбw�vk�Ѐ7�b�b�(�򂶵RYScH�Ϯ��	Q�p��#�zV|ZVܼ�;Z�`�+*�F�ɩ|�%Xd��;L�����ӵ(�! �vM}X���\��X��yJ�����u8���6-_��x��s���4�D����[��1'����hc��%�ធ���&�3d�sx�1�W̧�) Q~F�V���m�7����ϕ�_�d���_���z3N����v����q�s�-�V���d���g�+jڋ"ĕ���=h%� ��B�A����G��������HG��v�5yq�-7���B��r���9�I����)j�l&����	ξ�P/���C΁�sXP��ŖI��E��9��2�%'��`v7H_V�{ǅ�w�L�*�Ɣ�>�t�<K��g�uq��*nr8"}�~�{+\es12��T�I�8�����8���qI�Ut��#+�5�y�wv��k��0�O.�n���V��l�//.e�r�������r�$�Ɨ{�!��h��.{�G���r��?�]ޣ��9[�Ns�[�_����);�:,��j�4��T��~twy��ΐ?�a�r�t|t*��{<ud ���t���]�n����E Ua�_1	�C)ف�b��]�Y���n��XMw{��å��\��J�~����$S��eEf���9�S�ɗ�M���/�>�I^)#gI���=)p�]DRyV���sW�ĩ�q�IasZ���u.�Z��a��X���Ј���c|�b�O��K7*性��e�Ҿ,k�0䚥�|A�Ҙˍ�}�KU�t��m���C�KЭ)I�'�5W�}�s���9 ���=���[!`�7fA	����*�`l2��T-~<F�_Fh0���%#)�Ά�Å16v��w�������D�Ify�C~�1�JxR��I$T��	���<3zv�G��������ox,��{pPna����5p�υ���ur���AXK^ل4V8@��79�B�X�&^���_PV�ۥ�9;��&�Kc�'������S��Y��\����jc�*I0+3V��g�j��K�g��]8!B�E�	p�7�m��<Ί~zlɾ�5-�d	����O�YvM�>�f����靆�Ew��[ޭvܲ�-WbouZޕ�q���%� nWҬѽWW�������,I��w�Kw 9��=��[��2'�xbdϑ�������* ��� ����������U�c��IeKO�|BN <�4���q����L\��T����2�~����^8�q�.RV[�<���]`!E=� �N�_�$�[���,������	<���ht/`'���e������R[�1�-��o�"*�N�k��+���ٓp�D��M��ɕ�#�g����vY�VW�D�����Y���M�B�$��W����>w�a�(���T/@`���B�84gزeTΑ�K-��.ǃ=
��c�pT���vt\1���5�g]�������G\�� �}7(7���̅	�n���"�9��/��ik�/&!`Ӻ,���,v�����8ƍ�q�>C�'��Z��P�����J	�zG�?ˁ"�Ν�#��9-�-��R+�a.G�}3��2u8��9�b�_	[�p�8�H��-�[�C^���nX3+��9Q�O�o1G=w�J��[�F i����~���PB����8��F5�V~�:�b�t��Y���e��*+������Љ�Y���=^����`V�O	��+��X���
+�]$l�d�������� �� ���Ȝw;�pI�u�7U7�Hw��{�?�Q�ʬ[���/ex�����q�� W�vؽ��&<z�o���ۚv�[=�K]�]�@���Eӽ�_^�<��>T<w\b�@6HÍ/�I�V�F���KGW��6~�����hi�*	\��u���uM���Ž�;��4_�Km�XMz|�)[�[nN{���O���i+�/z^"a��~d��L���#ٺ�iC�}o�<�-�W�N��;8�}U�ÅS�����7�3(1�z#� -�����p$W��.�����H�AK��Mn�`��bO�4�1��ٿ�5������d������p�4s���Ɖ5��c��X{�Fi�cc{�:�B�{�fc���[ �p�,ꅘ�G��L�W��	~k7��|ςڿ�5~��~i��D��������Q��2q���mA�Y�Wl���ӳ]}���(�)���z���_W�p�IbJ���U���U�}q�U0/�n �K��O�/�e������zl6�n`	N �iE�03�@r.�Pd�+�b��í������e�5}�ajby��z��!�t|u�	0�+\�ѧ�~u��eV��i�3��ox��(=��V�o��Vצv�f�㯱Ʊ1���6qS���k�h�� �+\nmq�r3���/�d`������[���ڱ���B$���~��k�Bx��
Z��źZu�W3�r���σ�m?��Pj�=[;۝nv]{>[e����f;I��V��4b2g�U�`M���&�ľ[Dk�����d$�M-������A �\�����ѷe��证j$���^��gU�&� !�&���Dk�@��}D��ٞ�UبF��!�Ƨ����m��	�sL[��H��I��W��Y�����*EA�X*5�a��{��u�;aϋ3�|ˮ�&|��r��HD
�k�fp1M����4�,W泛��&)�Z��;nEn�,�­����	̺�I�6&S��	�gA�D+5������rL�mv��5�|Y�_{\��A�s���^�gG��h��}P�]�W8���Ջ�5�*��-��'���.��Z���s �S����Stt7�;A$#��&�u�G���[��}HT���(�!L�e/Z����H�_��{���%ԇ5N���W�IyI��)Z���O��J�b��>��������R�K������\Hn���z���G�}E�ihf	��	ש��="�p�Bu��B��]�pX]�y8v�/�A�@����X'�M^:Z�r��*f�T5�@f4��!�y����d(�LĢ`��a�k��b�+��%�+Q\DfT�e>.{?͂�
0ک��J���x����8�ؚ��3*cć[c��?�A*)�����a�������6���y�A����zE<i��U70!��I���!4�Hw��4��ݣ�;���;AGN�ֶ��M�ogg���X%955����g�(�x���0��q��冱8X�z��f��{r�>_��Ķ�1��y�m�`a�9��lH�8D[ϓ/mh{>�$�����ً���Lq^��ǒ�t��:��.�3�d�Ę?�K�YU����ԄҮ��'K�'�����-�5�D�}
�t�pC�'M�0@�"ڟ�U@\$~EĬυ��&W�b�����Zwor�_����a.{,�z���zmXJ��,��x�˂��cr{,�()��I����}��'���[
r�OCK?Re�~���w�N��-s�X�&�8z�h�~Gơt}x?�v�wYg=�z�u�"2���%;}D��l���~2[Re�`߷�RjWjk�8�FiP�+N��5i8P���]]t<%��z�&�3�P�]�4����׋=H�֘�hW�E�c�p�/��ċ��˼��%�+;��Rlۢ��CD6�T4�2XE��o����t'��bg�h�Xl����<��J:���o�S�CI�όJ�+=V�.���Bw�b�I,O�gr���,끫ID`۟��@)�걟͹��1�[��k�u�ہq��|u��|���A�A��W�L��T<��ٟY$�B�7�ᔔwDVzuYxqx�A���dalln ���d	�'����^�-j���޺ݤL��{Pb@n\��6�Q��+e*TI�Ӓ�H/�_)����Z��p�O�����?����܈�V���b7ĵtcW�Y��6�9�Oh�2=h�u�F�a,���I�K�cZ�c5����s�I����XD�5�bHٟK���	Q�b��PA�%lXY�tg��c�S~}� ES ���#Wd	S�if�ķ����gY��I��\�
}2S�R,������P"���F�(3����m=���"���ʋ����Vg�~�{�����j��ô��?����h�"%�������Ę#TqK3�K�C��B���q�so����p����v��,��Ĭ����?+hBK����>�Y(=V��MB0��g[��r�Z�P���8�L{��|�+�'��;�98���ߣ]�3 :,��7����2��*�ڍT�	F$.J��mJ5���gJ��zpaU�zs՜��\� w��M�֥���Y���kL%]Ms�?{/t�7�Z4�K%)/��,!��|B��~�y��p�)�F+%�6z�r$��y�X�ȫ�osd��"�l���7f�V+N<&����q�q>!������*��8���1-`Kx��y�&�{�)|�g�J��-Ye�[Q�L��;K��.=�����G��$�3������
�hV��n��-������+ss��-m�o�a4����v&F<ݘ��vۍ�ia{�U)��g�	,�>D��f�
e��gPdVSp6��_���K�� �����Jf���7��� ��6N:�Pe{j�
�/�B�>��p���~�KZw4''��R%����\)�W4'~���Z�.�}���E@�_����a�=��A�k�>c[�4-n��S�؋X���{�x���a��4��"�7g8
�L��ؐ M��B[��VB��#�^��b�5�s7\�U�c��B5gDh�\2l�V��<�U�p��7��� _����*����-�m�Fs31R��5?�:`_��.Г6!#�@������u��P��xNω��$�ʸ(�E
��г���eɓ!C�"q��z�V��q���A�F�����	����?��ݒZrx3fV�s� ����5R y�@�������x,�&����Q����	5���#�~�9Ot��2��_��ܘ&��_�YG���"}�'�k������_� ���19oOv��YX4/�98
�B��g���b5fϾ���:~��9r �qB����'1�]H��b�����XLL.�9.Ķ��g:z�����L��R�}������7��4~�h�Qi���[:+�#;l
�|��q�������2}���W�c*�~Fd��5X����N�#�B,��W���~��/�����P�.��<׊�a��;XeM��6��� ���XlW0 Ӫ6��U :5����gV#h4G�!R���lc$`aʾ ���ί�u?���K%Y'$���>S �	נ䳺`ᣞڎ�`-�w;�A��v ����F@H��f?='��׆�^�sꏕF ��p�e��N��]����lWИ6Yʤ��
�@<*��ῐ���޵O:�~WR!i�1Uv��WG������ŉ�z$�n����Bj����o����!����ڔ?\�ߴ�] c�2��O�P_䌏{����ϟ]��0���W�7�����I���څ*����!�!c]���7zhl�j���	��R�A*��~m���^*�a�+��>�ja(���X��NX>�N�xb��aA�`t�.bsz�:�"����^{��;vZM_1�Ç�$�vL�� )!�yc5}��W:��c�JM�k�����VV���27�t��,[I l�sr���q3�Ek�f\���Y�?�@"�2�T$�Hbig��=���.�L9�}@-LLe�DZ��^�#��O������Ո�w��v��2� �~�:B�-3�^���!�ԕ-���`3��C�N��"tAg�A�EVY�B��ҝy2~���\�K��㱗,�0{�}���iʻ���;���2b1���G�ҿ�ʹ�8�?H�r�GM��g���	�lP�  ��/�/z��2e�^��3�$gj�K�8-�N��2.����ђ�! �(��y��&ǞN�{��7�ק>���ݍњ��[�æ]|�_�tA�����A#]Ɛ[*w=,:^~H�G�A�gr����a*�űG�mZ�g~\��^��\�H,��4~e�w���rqȺ�Ե�ޱ��R�F�`��ɦ��-`�㭅����3�t��|��}B-t���G�I7p��
Vm9V��iaI��?� ͋���g��_5�����cn�1u?�����ňk��E���q���;@�e<S�_��O�Hh�U�ڔy:m�@/V�ߖ]�O����RD탣n$�J�Ԉ�u�J�YW	���=��6��Q��̈���e���\��=P��[c19���*��z҂� �:�m�ҧ�v, ���*�2�q]@:�va�F�K
��E|V��~-��F��i�ࡪ�x0R��ߊD�Ws�`�F�'T��|���������9�r��_�T�~����q,Q,r9G�����w��I>�G6���K�wGD2X].��ĳY����Xۜ���f�z��K��������!(?|S��x����oTR�"��~�,�߆�Y�{_�l��07��CQ֜�ќ3v[n8⫆d)W��1�m~n��;�������X�]@��8���m�{���x
!�|Z7zHsQe����o�14勃T�����F+Xح�v��>����Ԥ�"���c�i\�-�����y���ZIM�
�������_�UEG��	���Dڥc����3W��F Q�)nS�G�/���e"��m�tj�c`ﾮ-�~��%1�m
��o���r25�'y��9�~�S��\�$�KE� Rlc|��{S�Ŏ1�lًjĤ��X�ъ���N���1�]J8C����G)�=����ym���Q�0+��lϧ�+����9�Ɂ"Z=Y��8QpLR%����p����6�|��s��Y�������kr��L�Lrr+G߰��߽CB�2�W�/����_?����o����^�I0L)Zcuw�X|�?U����x�0j!-ꤐ��BOc����\~8��h)����~�_��&h;�b2�F^">�^&�,3XW�����,�+ݳ���ʺJ)�'����e�{z����C����P���t/K���Q��������~�:��
U寪��^E��c��4�l�P�;Xgs�����ְ�\�&?/�t��I`�t;>f���s4�cz3Br%wЬ������QV2c�$T�$�����NםCKM��x��ȫ�Mޫn����Rm���n�<�:X�@���/�L���r���Dkd\�hT�FB�p����"s�6 Z����}3Y��R��j�<Qـ�������ρxڨy�W�C�>+�E(l�\-��"�D"��k�Ir/�+E��}�	"3��M_�7P�ݔ1�	��	&Cz�߾$P��^�62z���xȵ��/D ͧo�d}�d�4�uyV>z&v�%3��:!��t�l͔ä���Td�sR)G�l[W���bF]:��O���Ў�L� 0Q��2�6ti���D �q�ُ.�������(�����Ŷ�XZ�L��aX�z�|AV㩲�4w�q�@��ƭ�l��¥}'��~��i���D'���A֟�i>��l��<��U��[��cK� �,�1؉;O��r���+�����0!�lOƇ���F�R���d�k�T?���jIEK���OC�a8�H�
6S���]�b(x[-Hx���Zl9�������D��t����-����ZjQ5͏�U�zjuOUr\i��1�H����U��/	��	u��ʿ��݅#��f{�J��dY����J ~qËuFT�.f4#K����C<t|,�� ������7� �h|��7|�q5>��%~��IX��j��e3��6#��0��+�2�`)��i���l��i���GL�Z��cV7�~.�!k\�B�X�4�����S�4����
D]�"Zfm������zڲ�4s?��L��9R*��=\+�{o�͍��NԈp���Á����4�rk:@�/�m�1+�8@Z�J���%:]��m��u%ݹ:�f�J���P,�g��w�����?��/8��
$��/�ВC*s�vI}ޯr��m)���J��w�a�e}.��=�?���(ܗL�4�� VZ���y�+oLH �76� y�jqzv6�?�e�y���"��ӂ4��ܭ��uɛeR�����ʅ�c�}T#{پ���'� Ӟ���H�)�T�}��B8��)�e�B�5�v��/�U48ca�6�ue����l��_N����F�n9d�t�K \�-8�:��lܤ��!c�G���p#�Un9���&�A
����j=�������� ���9�F�$����g�б)�}�]���(��7�m�^�p3ت����:�Q����3��Ǭ�r	8̒�J��dpfSV�ҲJv����/f�3^Y�rq2� 9�)��εÁj��ͨF�X�D�xg�x�^Ѣ!*5P���&��f�8A��JSȟc���h��y�*v~E+y�o�Nz�����z����QVg*�7��]�Ku��
��	giii�k��iv��7_"d�9Kq�+��Q<Ԟ�}]
Y'm`�S�X�llLj?&��lq!�%ߡv�F�ū��7�6����66��p�z�Wd�⺸�_�c�2F�61���C�����\��ѯ1pCg���q��]Lx�b�׊��y�RDR/qa��NI��]H# PV^k�7���Bb��,���t�����2Q�|}��Q�����5&���$j��R��4�x�h���.�^�"ۙ����DJ�?K��&>������7�,ٓ�h\Q9��"��b�&�i���|���)��<*esL?b��t�����M��t7�س�D]R"%^$�����u$[泐1w9���YcJJJZ��X�.��n���C�S*
J���᫩��I�u�U�����Wڢ;�����DX/�Fk�rat��n�g�z/��{�~�t�*>��NFf�"�.�����B�\�jZ�1l�#냳oT�_t��ĥ��j?� �vM^_���`�u�	E�H��n���u�i�=���X�0��E��9k�}���i�h�*?�3�#������s�L��x�N��U�<�>C(��U�eV�e3X�[a��O�b�Ⱥ��l��}h�q���l�����D��W�S
T���GվsS��]��+Qn��/�<�p�5�Y=�g
E��sM� ���vm�h0�)Zs�t\N��5�@��K_���kV��_�w{����X�}ץc���7V��cV�b7��2?���,����Wc(��*6�j��^5���C���6`�[����=`� |�	��z�D�}c�6�����ٖTLt�����]��<��Cm�Ƚ��ݟ�,��RL��b�doTc�C�i� J����b�(G(_-�p)���͑t#A�ߓ�W���s�Ϲ5�6�޺�E�����dm|{��E�U�.+��&4�3�\ �f�	����Ⱥ"O�P�%�:D��,u_����E��e�|��2Y�
]G)�7#�H�+�>k�= B�-�����gU��շ�BFm��kױ!`af�wsy�����9�poL(��K2��lݪ�c��M� I���؛Sꥇ���$��
�}��q��움]�b5�,Vd��O��)||%###^$w��;*v��cT=�(�4>P��hP�P�m[��h��Jv�>g����[��tq�Zi&���c�W-�iR���
�$ҽÖ��]�b�
�
�,������5(>OMAD��-�ck��qt�Z<��f��������.��O��By��8�A"�6�:)�?��w�>���wz��z�O������~"�d�J�u.��������'թ�n��谏`�qJw3���_�A��I�>�~�mBCH�ɽYEP�,Tr���]ѐI��>��7�ma��%�����<�d�z�_!lT��Sseh��͒��,l�h66>q�$V�f[�� o�nGm/qQ������]�tw�����
?�V�<��� ɕ����@/c^�q������P��t���z�k6W��9�?�oovC�CGϐ�Y�7�(�z�hL�W�h��&qy���=����=����>�6�,��_?Md���#Z!�S!����5�Nf˟�G��q�Ad�x�
>|�>���@/��o��/v��6��I��^��m�-��ԈVm�	q;Sn�o�e���K���d���4�X�~��#���)���]��#� �ˎ�8�Rko�9�W	�b���i�\cΓ����KY��~�N�D���c3��H���41k��y��P��NZ�r���!��m&×N�2��J����Dm����B�m)1�o/����3�^[��Ϩ�?$��?w��m̕@j��΂s�f��{k�U��n�M��y٪��X^�F,��'̸�0E�AW�~[�˱�LdM}�����5b�O6z �AJ7�V<nVS��5���K���������n���w��M~�|�o�˳&u������ժFX�@v*� �|δ2��Pwl@��X��y}�j�(�_F����+�$�
)���P��E���� �)د	^f��(d�zp���a"sJZ�;H@������%q� ^��~T�̴k��)�t+�uI��5A����smΨx=�Rl�(D�� :�1jU䡴��0I�
ko���Zu�<"�L%?xV9�z���7��B;�܋�P'I��جZ�����UZC�uEͨr�����Χ6���mkc���^A���c���6�sRo�=��mE^�HT�4\���͠@�G�?�ޢ���oV3p�����L�&dKK��aI��P��R���Y\d�Y+�W��D��LF��hy�`� {W����wq��1�%@sp`��黛�2��[��UwSpu2�s��.��/�9�,)yy��S�m���W���/��.�SZ)%��~P,�[G����d�5���!�ߍ����?�V+�_^�i'��y��Y�6��?�ߥJ �+�� �3�Yorp�!Ⴢb`��4纾�e�*/%K�kҏվ���ZӽY���O"�"o�F�9��B
�;��_Wԛ-�)�?���$RZ�.�n�4򷌌�,'w��B�E�/���/�B8��bͨO��H����$���(#>oln��Xw7�2�A�{�){�����5�2���gCnN��K������ ��� �3��h�u�*�Bdy̟�1�&����8[2"���`�稦����|b�f�²�ⶤj��i��j�ÙN��_:<f)��|PPЁ��L?i�׻�w�Dg(��fި�Y�?xT&��*x����fi��2�^?�
u�����0�_A�F]�q8��#E(lg)�����v��Ry��M�g���Ǔ��c���H���UPQ�B�u��0��ݎ ������dV)��;eQ^�S)|�g���[&Fk��u��us�ß��8O��b��D�]޽sx���o�Ҙ���j���2��/�-�ٿ����s$<�H����i�!����Ki�\ 
��}i�Ł%�@���Ë$�ۯ�����O7��L��*zw�O����ס��'q4D���$1ā����S�uj��s9F���Q?�g����+��}=Z�[MA*��WN$��0�Bm8�ex��P���W��ۖ^.0����<���X��g�Մ{SƆ�n�Z)�=a�c���Y������R���lh۠�:���[�ڃ�C*�i�!a�Fłr]�A%���R��oVX��x��/�>Y#/��~0�4�H_C���7�:����ٝ�$d!��..ˑ؛䁥��=<{��]��׫a��-�����>�o6s�5ro㬟�G��T�R���*K��G
J�h�;1Đ������"l���9�V������F�B�� Z-vG^������yI���7�GZ�Mx�7;���q
��I�+�`�P,L��J�4f(�?���b&���;.3���Ѯ��W��@φ����pg'�!}��m��ߍf`ApЕR\[X���mӝ���̈́_�n��@*���j�T��DK�!wk[�3:`���Jʮe�N${�p{dmg�q!�q��m�șo�!0J(�vx)3���4������[��l
.顨6���.1!�7I�V��R��8�9�_��M_jjͷ��?��3����{oѓH-z���#A���E�DD���^G�ޢ������{}g�������>g���>{��hM}�nY�0酜�� ��Q��������eK����6��G���	���K
���Q��#���Ir�'�7��?+��`C��c*�}���ԟxz� v4g�KE�&���k��q���UW��q�{���_�ld���w�%2�p�S�>��{X�xA:Mڛ���2V\�]�ꖕ�{0	<1y��o�yz������	Q���6F��r}����u�8Ib���b��م�����9�Y��0_>�鿪��*h}��lh��
v՝���{�a�حƃ�J��8lsL� �A�W�H�8�LM(�F���$�����J�`MQhN*�����ɉkso��RS_/��9ѹ+w���5�����K񼽪�C���_��_��[�P�e'�e�餳�f�����LD{�\o������Ǉ����V3��Z�H�o�>��ײQ!ڶA)<` �ŏ��ɶ��e.�����ן���D���IvK֋��p�ɑ�x)A�/�Zin���m�'ci2����S<��ñ���z��MS>�#q���#ҝEz�p��[���y�r�`�"/dL�8�N���,����n/�t�ղc�/K��zP�����o%��:��x�j�%؍� �V�̠a"��;��K]T7�Aᦱ�;b������P������dY'-L�w�@[:&�����&%��+�V�fZ�'�?�J�z��ٳrM��[���){�Lju|/����K�3\���Nd����R��|�1
��a"�z׀�J ��Ճs"K`m�2���G}���_�䴡ɔX7�*����������������h\����qR �)�/�p�|;r�o��tص�e�ӱɃ����֛�}S���JFi����w�����<?M���-�X�H&]�b棉�.��͐�>���Z.�)�VU�z�N����$�MA��bykC�!���@xN!��E���f�9���4�҂z�rJK����1������;H�e|��&�/�E�ȏ��:��ೳO�<i��ߨ����ӣ<::z]C�C�TPP�<ۥ/.)Y�9;;yw{u�,�E�,���J���#x9R�UY�R�&A�����&<{Ϧ��~G�4�:��J(��ۡi]����0�_Z������|�_��;W�6-���x,�8�8�T����w١׫m915�o2��5o(��F!'%�˼4�A��9�h�q�3^��)횭pt�턲�ؘ�D�����ls��QNlu���!��$D ��k������ ���6ʒ...����[��=N--�Q*3y�� ^���Da!���(ZR�y~͉z�?\@(~���^�fg'��{/TBb�	+�B�*Vf�p?4�ef`�w� ����n�g�ms��g=J�sx|�GDJ����ʿ�ޚ��-���8���%3[�ɯ종�����{$%$F����y���x����y�I��B5�_y/�F����`pBb������~O��^�/t��+�u�10D��奲��i�����^	�9�3$����hu8XW��S��j��X_s6E󇗻w�F�G���kdX���"'N&7�(�׸�n#�$>s�� ,;���|;@c
'٢����`s8s-��gr�3���^N�Bܾ���~L����k�:Ȼ�k�:C�*�Tɩ�6M�}�<ݍ�	�9����11�h���6�|��SMъ3.RM,�$,8rd�F]��6:@`q�b�����n)�*�8�6<�+Y�7u�7u��я�U���g}䎈�.Dsd�O7e��/ ��3����4��mz�m����߸�^������{ ��Zh�|K�u(ޗ˔�J�� E�$)�(��ǵ�Pg���ǿ4�����n��NHBW�=,��k�����Q��T~g����r5Vr#uKR��3?"N�ʶ+j�氧ɨ1*!>���x*>U��jgdW�}�����J�r}�,ٚaV#"j�{Je>{~<;1�jA��H�b.�<Uf�Fn`b�(���\);��2���6��K^K+�y�De4ۏ;V�|���8���9F�4���ϣ�	ƧD�>�*}��S+]3����~mu���ĕP��\�����󾤤���­NmzBB*���F�b�݁�ZZZ��E�s���?�v�B�b����7����yF�B��T����D�M^�	t)
�t�E�.
˰��+"nϾb�2����`�7��K�;S�!X�}����0\���u�{aZg�{tɸi���]�x�}c�wXi�����@c��ø�'C��*󋺃/ͺ�����5x{�	`�H�<id���7�pm���KeTB6
�#֡�6��;l�b���[��H�Jy����&��.���š��''W���> ��k���#~�q.�=̬�U�Q���[m�9��=��'~Y���[��k��D��*�^д�qՊ����e��
Z�3xun�2]i��������S�X��|�w�_��o	��a\�DX�X�%$�n��M�*M��.�ɷ��V���ř�ô.L"�F�	i����x�Z�1���V�m��떇�~r�
O�-I��!&��w�^��={g��=�������#��f���QVW~iB[�;����V-�kg�:靿UL%���AV<�P�_����rs[�a��G)�~����V ��mp�Lq
��ފ��v����N�w��K�t����U.���u~�wH����dSq����,5[=W�hM	�[�������mO � �Q_R�_�@�gs�w]��ԃf#�sw����J������f/15<�?�.&�uc}y�.�� ��NqI~��0�P�c����ٞ��2�S�G� h�AD̊�N�;`������mvC�$������g�˔����|L���D8w������;��b�diGH�N����*�\��K,ܴo:H�ј�^;3���6h��K�g
�C?��u�֨`cUz�jH/��W�oV��+q�A��*�s�tp�TQL#j2�D���̺VfD�B��k�<������W
 ~W�����.1I�T|���F<z�yMb���	�y~ն�C'��뫊�����s/���S����IB�]0�;[8q<��q�FGE��-� �ڽ��
�HL3酩aS]�Y�WߟvA~�6[QZ0�-EO�ƍ��s�c�T�"����s�uT�����)<��'BXm��6����f83.�	�Em`�j�h6�3�c�˭�����_F��/�z���vgy#�	˳ù�_�{�B��/����Y.ꤟe=�	28�=��貓��`�T� ��~��&JT˨`3H�}u�;��η��Q�E��@�zv>�4

S�NK~��Ws`�b���1��ҹ;(���#г�8�$�|�e�0y����&�*�|�'��G4�q��:�Vi=����I.7���/�qŶ	ևZib&����OV<A<w��)t��Y��[_���FD���yH8x}�4BDR�S";P�"n��;���G��X�!��(�:�3͕�(��o���&O'4`O� �;�^s8����uv$l�:�Ď��D�gy�v�����"رԅ�Y�W�i�`���1�����B��|�͟��|��FU�kjz'�^c]T����w�\���?�:�||����k\e
��}�(����T��뇽c�7V�վxϣUU�m�L�x���`Lpv���U_q 7�6b��W�����_<��	)��[�u�����п�-�������{1O��A^�����O�Ž=u��#��?��Q�Q��R�x&ɄZ:��+�Lsh��L�\Z�'��7���Ik|�U���)ڣ�ذ���f��$�^��i21g��Z'�#��������׀���>W�s�7km�A��ѡ�8R�O�D�o7�bv>bk&=A�|I��"�<�m �u&0�랡�o��nu����:�f�KZ��xEX���{��
Q��a�m����C�-�t;�e=EV��B��/Q�ᔐ��8^��g��Sşp^�މ��t�����R�bO�t�ssv��!	{�Z'Y����06jc�q;��.��Aeo����w�d��k���.�:�[�Cm�3�Q	}����-m2ch�n��߶��%�\��?F&~��L>|\�����f��[����3�+"�����(Z��_��Ŏ�	�=M1b�\�/^�(�u����R�2�YvnK�|+�g�T��n�B$��x��H&g����h% h`��D��ﶷNN,�"���`?-��N�b���y-�t�.,��s��}��H`�%����&��ٮ�3��?e�_��͒B< �}7�����; �g&qN	�b�G0��=m	��Y�������q֨�~ei�7bIE9k���'k�F�������P➳���Ew��HD��j&Kxx� ��2ݚ�8�/{��5#A�߰�y+]���y���I��3�}��/�l��F�� �$D�O~���W���J��%�&�?H��Ox���I7��,��+NɿJ� �#Kd�����D�����*j����d��rE��A��	�Z/�}��H0Z#P��3,>��7��DK����_r��,���9�d�L�p��X]_�J�i�ãP<�q\��s�~��S�m)\��Yij:�}rIPyDр�f�����S����{�2�S�$�NZ�Qڡg@@�"/�Ct]�d��t�V5�Gڜ)�i��Հ� Zw��n�z�����q*=3.P-��\���`��W=���,o}�`�6���������"*�_s'�t�2"�y:4�b6r�ik��Ͱ��S!�Ѐ��	�ah屵���Q�cQ���4���]G���!��	�\�%�Q���p�O�J��?/�'�-S�vuay9�*��6<҇�n���!	�d�������9w�&�wJO|Y�$�bw�a�(�y��H-�����|bp7s����@����*X���R{������Y~y6>zĚ Vǳ����F������Y�ɿ� =�(���Qg\�m��Q!+�xDb5v���x��^ ��J��&���j �jqK�fSƿ��yC3(�؁8�Jz6�̕et�_s;���"�7!�uT��C�!6�~�{1��j�H1�����[��;`탬7t?~�>�z8�aq�{u�7� �o�����Õ�f!T�Q��_�R$�<�*�u�z�W����/�N���)��z������Y��&���M��X��3�P�">��0e]�+���00�����M������6/ND�����B%��h��I�d��`��µw�C����s9��X5�B�Z����~7���?����6.`����_��"�1���n�6~�����\�Ĩ�&$�?�U�M����Nj��CAf)�%��r�z{��0��%��ׄt�2���I3.,,EJe56�P��At-��F��4�&gg<����Ʒ���²�EΧ�I��<� �(h�	��$k�sB�)�=$~#���0���7�9�/�q,+�c9��ʹ�U�.��/��E�S��0�P4wa���n��mFU�m�b�>9n�ց���ި�@a�����(�P�X�l9��JQ�B�2WJ&�������L�H�>�ϐ��]F-�9�{�ɾVR�?:>�w���s� ���r!�|:�aS����d��s�rR���S��I�Q_�L�yc�)M��i��n�6f#iqȘ��ܙ�bO_���2�����ȟy�8��V������s��fۤ^�|��Q_����*3�
۳��8���6#�Gl�Q��t�����ŧʋ�:�:�@\(��RS_�s�%+S0�+Z�B-�Z-�d�b���\#eggg%�o�[O�ߖ��&�LG��$A�G����P䯞mb���23GJ�*K�ﶟ2�l7���	qq7r�Q�[��mMz�~ �?�J���W[�"�X1rL��6%㰔V�n�����c3�=!V�����t�(��.�T�P����uض,�D��6�a,H2� �������vG7t�ƒ�M���ݙ���ȨH�5�v	ʝ0���zT7D�a�K��L�SpGQ>�D�eJ������ ��(�p��1e�9�>��b�N�N�z�N������I!�3c�/zb�<������V��VPٞ2�������b�����5�k����@d_<���N��^GlƿvHRB���#E�Nr��:E	�$�ϟsw�iDO�kp�A�L��±�'W敮����֘�=��;���jHNN-�d���D.�j<e`B�8��ۡ<g����>�/���V�a�q�
��}����FF��O���A�^T��{��Xg�'��#Z�}+��|E�m7�ݧVkE(�YG�2S���'7�SC�.S��j%��^�u�[��<��;MJ��A��rr["�Q�u&	 ��G�;��|�;'���s��Ѥ�E��D�����Y��؏�w��O��o����g�G�֢m�D����W(x=���o�e�JӊǙ�������A+}_s�4G�ʁ��D��OH�JɋBŐ����M�x3{��*��}ʇ�b]36�Y�D�C稼OTm�-\]u�
9J1ҞK�����=��l�����ޟk��O��G�}b21�#d��Ɵ�R����KO�o
������Q�m-�����M9/��l�|:P��ނ��݃?<��q�VB�RPT|��>���~۟u <�"����ayE�n��2�G�~�7U�^b��p�s����xr�E�sw8	�����?��ԉ���_F1�����T^ؙNT����^���:�j�p�l*A��o���;pK��("�ݍ�w��i?x3��F4brfU���0�1�ƈ�o�ؒ�� �*Ҭ�b*��Rp�03{�k0={z���%WA󆳺��톂��L�����Ǭ�h�i�Cj�H�M�fǩ��$�t�l�lϐ��ypu�=��d$�ӱ������5�x��Z�4���8���4���AZ��dlޯ�%���Վ%{��&R?��U��o���x�B�)�@(8~T��
����'+}�P��� �AVzZ(�,���_�A!Yx*A��]��d%̹SvOP�[��A�x��k�O�)���@�pLL���LS�u���W�6��im���������G��C &��9���YE}/]�o.$BAj4E�y�Q	�6�2U7-�a�sk�2R��P��fIYV���EW ����wzQЛ�����6����i�䯏��&�D��֩'d��
ˣ�F�P�#W�Zɦ���'Ϗ��y��rG�@0^"RR�XN]ug;����-�.:E��'x6��Bg���{P	����V�y���=���]�k�~�i���Aibrk'��1:n&ߧ��YS�):ByYg�҇�?[=l�A��"�5���!0k
�{�����o��H�[qiq������ɷɩBڃ!������.�.���R�u�X���
�:�f�ĢQl
�� ��Q:��\��[	H�Z�����}	��趤|�P<!�/R+$G�czT�j�>JIύ�B����@�dI�.�ܦ�&���xkC1rw߽]-���]�4Aġ܊��|Yv�0����y֩NX��b*�`��<�x��	��>~�ɧB����$,*�r�܉����ú��ۗ8��O�ASL��s����Z}1k�F���t�ǿw�~KD��t���,nU�[-�c�Iԕ���G�|w7��I�+J���i#�&��5JH�5s��?4���nJQt��uqq����9�T��Nf��C��Ӳ?r/D>�V-�E�Ț%��d�N�3�C�� A��~��yFp�A��9��>f�,kEC.^xA����S�ݩ�&�0�i{�r\�x���ZX���) ��Y�!<�1=	A�s������^)f��u�Y2�K�p��Z�bl�������gB-�sr����!Q{Я^��ޫ?�P�L�'�[;�v��1>P�ѣl��л��Q�αv`���&���7؉���˱�{¶L=�r���zG�ϟ??�?W78��7�<�$����	�gY�\�qss�]ិW�Z��C�E앒��������F�ɣ/����,أ�G��t�Q� ��9i
V���\����C1��A^�k�$s�	QN���,n�Aq"ߖOEc� �k�1w'�@�
ӓ��d� �x�A<��mu=Z��ˈ�A�����:uvO��B��hZ?�:ԝ����m�Bg��;�}̄ǒ�Y{p�S�W6��:���N����4�ߢ>[���QbX�45�KXOZr;M���.U(.VT��K.�z�/t�0�`�@mO$����i�P]Z%��YM����6vQ�te�[e��)!�j+��O��gE��uII��]�/f�=]���9%!&�@9�Z�\͉>��*J!J�za����m(]�r���2B(yG?��c���6V^H��GBˤ(��yp����J���h�/��K�
Ry�!�5�Pv�tb>�R�O�YP��+�qm�,�!��Q�ns��/��I�:��K�n����;�O��~��7�̞m�B,A��"�}GPIU����8�@x^�o!�M�2���2r&&���('���Ŷ��R��'$t2��n����Q�8�i5��B9�)�i��@��(���+7���h�y\JHNOO�@�iT���9�`�\�\�/jӡo("��~�����k��2�����;�o��^?��8�A1�� �hv���w�vr��L��أr��_Rf)Tfv��"����]aP|������@ ��>���y�6��q�5E����[J��z0����o�z��H�/k�cG�P*�cN�p���ÏF�2{�0���5*����z���x��8!�O����xpᅻ&���3...J ϲ���>O�16xB8F�lO{��;$���o�#f�����ΨSk���.��Oz,R����������n�u�;�y����(3�-,@�bY�؏陙{ �:iF_�
��kQ&�E �X�ޛ�n�3�<�IR��"f�i�^���}�V��_��e�(�ZJ�	}Fʕ(�ѥ]�q���A�Z
���˸��QZ'Պ����7*�����l
. #�CAx���H���}�`W]�G�����O�
���ԝK����ҹ&��� �NO�'^�}��x4Y�n�B�syP����ҌVηF�=�q��ۛ�ڦ8�ߛ����l��_tL�F�L2��_n�����5?��`������4C��E-��y���l�껐u@�zt�r�O�b��F�i���Y� �����F�3-7{Z�����\	f���U��pv�_|,
�y�g�<�B~O���q����uH%x���\�Ȧ���*�ל�ڐ��Lby��U������k >%'o4"onz`�n5[;_�n^�0�L�uyyt�8���ߛ�����=IpR�j�K�(�ʮ������!25��R򍅩���h�>d����1i5R&�ht����7��7l�ZG�'�S���pjg,%h�8ǰ��6+	������ag����V�9;p�Y��Ly��,�����ݓ����,�Y�#�a`d<<ZS��	��P6�nL�e�e}L�>#�Û���p3G~G���Q�*6��+0�2(�D3�i����F�0�<k��<y�,�$� �X�呣�j�#�"���ޫ_j�T���K_�#p/6�ŻM �{n�݁{X#$����?�ﱏ^9:�Ⱥ+��r?��OD�ٟ������=��I��8dؖ�ާ?<7���>K]
�۝���z��7Ω�f�2�\{]��YK�c�� ��i���A¶y>L�ub�%�M�1VQnh��.Щ�DW������R��g&��-���>�z��5K$����qa���FIF�����j�_�<Jc��,�aN/���p���1��E��~O�a\3hO��D*��J�[��t6���>��L��V���p֚��Q���g��lR������X���]�m-����c�j�3���lw&x��nP����I���Ѫ�?�����_�u���k;�(%Y�����sbs�7r8Q���t ��P��B�զ���c<t���PҪ�ož�*,N����)����n��`�A�*���%)���3�)*KVr�E�h��W�\�=bz�h㽥��!HK��3���%��@)
1�u�wWz[E
X�L���8�&Ys#�1%uT���Z�˞��-G�5��|�5+�k�7�=#O�V�5«+_+�Szn����t�$WnG�<��Ep��V��D�;�T������7�3��U��J�C;ִ�/B��{@�����ܢ�vL���0�S���u�^�%}h@i�Tpy�S(
���$������
E�Ũ/��<- SR����f�qK)j/����/�T��Y���+*#�0��C��0e}ߴWs4u�(�s�&��B���Ɗ�єV;s��ot]l��(f�����z_m�-T�3]e���B�B�,�	7j�@��̀3**.����@��`d����� ����2.�Mǰ���>��6(�=�1Y�5!y:;�O>8�P~K������k��Q��@v����T��9���^%�z�-��4xY%��:� ��c<��ᑛ46��!c�;*�V���[��J���7>��ދ�ܿ��2w���h���u��7EGfS�IU�,���	u�t��?[8��<�b�zs���Z��p?~Y�jc#37/s�&ݘK�����ڴ"OZ<���C��q%�6x§s���5���{�
+��qI'�凞TVLD�'"b�nGF���g���\(�1X�Q�p�����,hS(���u�Л�P�*���[Z�hm}�CU@��-�^�Dڮ��ݓȋl��ǘreؤ"@���Y�r�������gi����.�(����}�G03����S��A���)t}�#��\��N}$����qd��5sz\[�����K	���Y�~�dU3b^G�� ���{?^]W�X�3���x����b@�;�k��J��&d@+F��$�#���&�C���� _�@�0u��8"P��ٷ�?���'�*�#`#��L&��	�ΪA6J�9� H�ğX��2���MYږvO$B�Y�'2�.C�;��Q:Uܣ���?pFm�d�h��ɗ��\���X�o�����p�!"��&Xwn�����&˹�Y%�0�`��)G9!X�h��C�[���_L�R�,�Гף��n}S'I��(�D�P�e�M[��]�e��:�5�����`R%D�cgVN�������Y{-pr��<�WC��sd?2�E���H�l�'���w�����c��:��^��fӺ1����y���p-9ߔd���D�z5�7�jQ&//V▩Ǧf��|U��9��Ƚ4`�ӗ�b����[o�S�������M����-s�[,WX����$��1\�!sz?��\�؅�Q�ϟw��"S���[
��u�9f��<g�8	��8r��r�ݖm�D����J�,b��%�+�v�8_Ё�}ű�ߓ���Н��Z�N��h�"*0:���ھ@�!�7�$;�:ǅ�H|c$�����r\����?��A���4N�E�&}nh�V7�>f���Z�̗L��� �C� 
�芧�FȪ�X�����c���'>���~��4~����M�X����#	p�c3õ���w���p%#Ƕ"7M�ьR������͐��x��j�]h}*��a4����l��P�}	�U/[����xS���12}��_�=��d��˧����1[�l.�5^+}�2�Q;�Ȅ��vl����:��׿�w�qϨ�z����ͪ�,�������;���X~K���T�R"l�_�OÓ�o�L���m_��9��b�v\�L�5�ҩ(� A�a���FU�{����\��O�N�=��p4&t�kK��N�%��Z!B��&VP�����tx��"�,��|���ʼ�m]�+��7�:�@�����C���u�oR��PvOZ����+� ��(��F���"U
� 8�)8/w� n��:lZ��	��VwJ�Mu��tY�mf�o���"�:I5]?�p-���H�E��g���eyK;S�w�x�SN�����^9���~���Go��A���b�����>zm����I0Y ���冿�H2%���M*�Ŏ���G����(�lOk���?`��"fu�8\�E��w?��t��c,�}w��A`�&1�&���\�~�G�r/����H�4!f t�4�H˒R��}@&q����ݎ�.�C�<f�ߕ])���(|1�	�1�$���8��2mq�s�}S��5F�J����V �U��m�����?��~oetmm������� �60��I�9'Z`\`����{κ"��{~���[��N�S��[ y����yI��U��!stK�����#)���Y�$��)�(.� ���%��*dF�\���2��'Ŧ��o�޿�0���!H-&��dڋ��Z]���`$J��_8��22�tiL�T|��_�_������ݥ��7�,n�o�Ϣ�� c�� ���ȸ�����'䖎�+Wq�A��}씰��?T�%^V�E���Vi8�w���ʠ${����]� �Tq-k��6{��1Kf(o���jOk�aaM��Hy͛m%���T�7�Ӻ�[pGa�����b�8G���}�o��XX�|�ú�+c�+�Bfy�>��N1��5O�,e<�%��hn��^7]�8z��x�2� [���x���T���oy.�K�|y4������Ϙ�.��]b-W�S� %]�do�g9V�{����N1�����Q2|e��3o������%� �7BXs	s~D�vy`��^���إ�Ҳ�e��ܘ3�{F�>���/��>=Yߜ%y����%=��Z �ƌ�=&����I�ܽ4����[����(��#'N3ÖK��ѣ���r��?�!���O��3�6̘2"�Cep��/�I	x�qvGv&�����K�犜��Z�� A�����^R析��t2�l��]�f�݇W���Y�{z���*�>YA�jΏ�~�V�o�lk5ӸO@�m�&���~k��g��/��f�SU�[aC=�~�o�'����k_��,�0UiҞv�o
�%e{�-b���W�k9E0��l7�9H���E�o��dR7�Z�@��9����w���(�&)�ft��P�����'���Fe�N�<i������1l��*D��MM��W�,�Nx33^d�4 ��[�6l[�l���ħdsqL��w~���f����'Wo��苆Z�N�&��,���$PH��^��ͻ�<���Ր���/#�R�0#����X�G9�ԫW�m�ug�4r0C�y[O��F4����4�9s�%�,����2Vh��I�t�����:�A���[_q�y����Gd:w?yG� >gA�d��v�Cw��! G�	<'U��:J�/Ѓ&)q�Ò�l|Y��mV6��T���~���yt��y������
	E�`└��Sb�FS-��T0g�M`���c�c��&���v�w.��,����b���̴�.�Ż<�_��S�`�?�C��k.A��Ϟ��
��B	��cIᘙ-��.��Zy	¹�f$����}�=��e��[����Ãe��÷UUU�����7���!242J��lq�hn�Ӻ���ly�`�9�?�a����y��筨�����"��b�����90�����J��[�7��������[1������y��@Rn�*��0�(|�z�/�i��LE�&�h_m�O�>:j�h6W�3=3}{Gǃ��Tn\�Sޤ����u����9����u�9|�|qd�|4�Z�!��z�[�=�y�kr�[���]ћT�?ۆ�����;��B���5��JI �d�
�=�7m�C&�!����＼�g>�揿�I$5Rb�/�y�����u���'o�!�n��q�|A�r��	o_�☲`n�880{[�'�o)+#��<��o�_�Ei	G;���n��}_i��q%x������ԃ��_v�x|y���G��K��Y�V$�f|�[��Q�u����v��ʔ�Ge����_�DCK���c��ż$���jlj�éc��H}���Я�׫����{����o=��yX��X(��{]\[]<F�w������SG����F*6�܋��[�~8CC/*QLW��m_aʥx�o�Bg!x����"?�����SR�H�oRgG������K����,�e��/*���;L����F����ˑ%���)K�<*���R�o�>��j��lo�V���Io��IYt�xp%f�ڴ '{#�%�"d��#JE-�5Jv܇\C�8y� ������D$�9y-��|J�����D�OG$E��n.�J���VzY��67mm5��6��SS;GG�&���]��.���1P� ����K%5�P�g���yg��QW'RS_o����R^Z�ty�1��Z�x�)�@��P������.��8A9 ����wB3�xg���A�|ځ �p��W���Ʊr��֮�Q�瞔�5�ߚ&�h9�!�E=P���vg�~_8]~�3�Ǽ23Q�y���n�!�ڧ1���y����$:&&�=C#�{���
�&�6�_G��>&l�M����{�p5=����v�j��z�[�g�&��Q�wr�(���aPe�����b�%܋!�T�KQO�0G�Ƥ�`���^v�Q��;G.C�c�y_��na��3<=g{�������TS=�444j�k"��PY�B�¬�p�����:��{�T9���p�o&-_?
�O��֖�I��k����o��˟��1?-H��1�ܷ�ߍ�2N����l��^��������%$V[DSK�d����|���"έI�9�?��Ӣ�iZ��W�E4�?+��'p3�y�[4�N�����»0J�j*����ɔ�O��{�z�I.T_Gcch�e�Z:7�v 5q�MGs#Ύ��DWـ�_eA5�z�7�f����Wv�%�8�(
�ׂ���t#�v4|}��(?(p���XA�-���>8]��ޜ�����>kY|M��m�<m��#m$���4�{�,^Y�̔��eE�sg��p�ͯ���{�����V#�sI7��7,�S'���Lہ΋��4��_e+/���H��_]�t�9�K�<g?+%|��\����Ua`1<ʯ
p0��9ğ�y�;��ʩO�*tǛ<88辣�8��;X�L4v��z��n��q�~v�K»i�C���$Zv�RS��P{rޏ]Yڿ[_D������'���[H�D��Q���G}���es����=z����676��2�fAߞ~�;�����!11ۼ��{�G������ȑ������:G�h㤠�!C�N6��W�^d|��֎���r{�//�܁555��ՁD��0�
���P��H
G��pi�pm��m�Rs�-��#QQ�bi��0�g������v���}�⠼�L��Y�-)�́��X�:N��ꣾe���*@�Q�'	�t)y:m�Zdü	m;�J)�b��U��g�jȪ��*��)W���-���?ƅ�� #Ejs�gz��j�����6�2��.���|�����G�B�p3�˭7�|��������//-$��`�"�u��|�)�n�,�]ˍ���G�PG�9�,��X;&���|݌�<ވ���2����ν��0L�R�2OW#& �ss���j`oَ��/��e��_:[��.��i%�z����������-��n����{\�ܭx��˸�G�ߪ�5�T���gf�����#c�Zh��z��S��keg׏v�U���]1%����>0W�ӗ�s���`5�j�*9�Ih)��^�[��|RdZG@���	��j��ׇ`���5&g~��^��[��u��X+��6�.D`�j�NlM4��6����H�O��P4�I0�+�a�.)TX�{22E���ھ�8��,sNJoI�,�W�|�w>� o}�X��i�Wo�+|i��H��k��5����!�<?�0��ͧr0 �d�e�06��	w:0@EM5�������|:p<��〮2�09������4 �[��B��P��V�ǝ���@��]�紿��|fKۓ%E���J�|oFH^35P ��=�iqC�H�G����ސ�VJ�;�l
v�8?(	��k^��<���s�,U;���8����S����HZ�?k'I<��檅��~OzoN���
��%I��3h�qO]:|ll�B2��H�����fpa#��w�y���"9)��&�4%+,��x�t�lxU�ҹi�8���	җ#��C��Ȣ���]n`z(��?�mo�	ò�£*�	�P�+!DVU̓�����'a�$�±����"�bn�L���y����_�.�u�e��ޓyΆԅC�_��M)$��h���u^�!.��!0qM���LF�0�� �TS�)�z�sű5�Y�D�{�����F�k'�i�X���_��xć 6��rź/2�#m��쮞�a�!!}ǡ��M��ݪ�-��TH��Z��;�P+؈_���䶋�8Q��#�8QQ��ُ΁?a	b5�_��e	H6.��?u�ם#�Sp:n��u
�yo�ݻ����*8��E)HP������)�-����+�q��"��ri�����M&�ZC}vQһ��e�?�����S�Y�w�O|������?BN�O�Q��¹�$]Jٵ�f�/˥�����9��+s֕g���G�u�C���J([ȦP���EHFF8;��l���PvI%�y�93�Ȏㆽ��-�������p���y������~�^�.0�7��N7�t�TE����8��?�Yp��ޝ����~�IL��'���wg�ݛ/�Th܃邟�"}<��N��Ê_�M�b�H��\��m$Dw&N�>���t!�7Bk��G�]s�zo����DQw��D;tO�+�5$T�A��/�ۏw;���
�{n�k�.���!<b�m�584� �c9�) '�l���
K�����<*�k{<㩙c&X7@[N�8%w�5n���vi0���:�����C���oF��I�S�3=��{�+j�=��OD����t90���qp+m�X~��lA"���:�y��ݙ�!�sF��_*u{8��gu�*]W� aY�7|V�u�"�S7��CL���^�Q�O�>���,�~�'ާ��dgm�3�+�fVV�}.���O�);YӉ'ȿɀ3�;�wr�md	�̷cy$6���(��~oj�&���Ϙ8���|��.)kOK�m]�$KH2�Һ�nv.���i#���%��fb����srU$�i�R3o��~!��7���P�K�y�d��U�:zs���~���/R��v���:�X�A2�B�ٹ 2]">6��ٌ&bd|+W%�Jbbbq�˳ Kl@�T�{
�%ꅆ�Ʒ�P���_��`�*b�[?���(EQ1qm��[���R*�a-�~���<[&3qa�q�9H��m������s���;V �N��fu=��=o��3��%����1�ئh��LȊ�VB�b��I5�:�${(�*�{�ݫ��N$θ�q��+S�@���n�㌑Q�������j�/Z@��|.1,���.����-�y�F�3�H�����������mCE����dM�yܴ��7���Z�]�D<?��M��Z����e�JN�u��>6��(�ǻ��6ҊJ���Uq�g��oS���bb$��Q�]Vv��^OZJ*�7KB^bb8��}�e�3����ܣˑg^���SԤ39{��ki�o�_9B�B��8^>�j3淍2n�{����N��������m�Ý��t ���>�QB����_׆���SWpo^x�d�5fl� �"����#�̞_zd���&�;�Ւ�j@^ �9���ύ׀Y���"����򮠠�$������YV���W+�R����_��TUk>{�K�3z�U0�`�ڧ��6�f~�a�˾A$�W)��\T=������U���'�jc'L���]7V�A���}� ��%ր����`!V�h[���_�dq���Fɜ���z�r'��B�R�4�>�
��W3�1p#?�\W���rX��8h���P&�?��^K�����~�K?�7h|����D�nd�8��?e�cOR0#��2�����k�B�+�G{�uc���CJJI��	������������Z��>x�e�Qڕ��g�SOa��X6J���;����K,�9<���ҍ�߈b�x�������'(��ƷŁD���������T�mD��>){[�L����������w��{��&�F�/��R�;ż�iu�k�&����߉%;�w�siǮ�^�}Y��޹�}K+\��T2J ��IsU0ݴ9}v���e�fO����T��3+��Q=��X�0�2��5.� 6��Y�ҸM��q+� 7�*o�T���<Q�+�;e����`��?u��?L0�v�ػI��b�zy�dqu��C�%�.��>�/	=~'�T�6x[ǐKB�KU��Sv����[�q)�nzo����K|��m�8����R�`�̔��:` 1��I� V>�P�ȥ���:�| �d���Q1Z�2�u�2T�,99�,�-��l`��t*�"���t��~r���V��D���?Y2�:�^3��q��aQ]�I�Uy�?�F�{q���wl-�_s>:��V�_u����ڗ�0-�gϤ�u\&�(q87���R�H�rv~dd�?D�WJ�D�I~��΂�O� h�>�T�$uU�6�x�	/���� G-U��$�R~��z����<e����򹌆�
Z�'�n7�b5޿x�ٰS�@@��&m(AH�r [�{�� �3�9E!����B�E�_�1�wޑ���Β+r�8��`}tR7��͐v���`�o��Ԁ��t���G����tRi�8�#�(����t��ژ�J��')��.���:�
qzwy!q9z?o��C���O��'������D9�������>�����r�����T��Df�G:���s鹒ᱺ̱�Ci.���=H����xT^4�����,s..���-�k[%7�Vs��џ��L��ߕ�� �������t����6��HN��T��$�V�v�]o�ǡEX�#�R�]/0��GKMET�CV8�^�)|���|X��^�����xA��~G֣D�&� �.p��t	_�f؂��WVA�^���Є+�K�ܖU�i;^ի�1QSS_��P���#^��
e�_�jh�W0������l�z�`�h,+N'QV���V���';�n0����l
��~�f��V�#+r��3i�g��m�_�?L(��T�`�]t�j|/K�����z����r�Y���eF��f�l�gJ(����6�;;'gs��[�W;	4.�[7D�6�|���X����8zI�AȐ^���qo�N#���ys�ٞ�MT�퓿�x�C�xi@��ôz޽����ф��Q�X�Yէ�<J����F�?�����*�����j��W����Qɏj@O�p�
�	�\}1f��Q8�Q�r��ǩ���דy�)o�C�-�3�u��A�U��ؑRWO�e����č_�>��M�Pz�-w���ޕR��N�Z����Q�^�x�Xkֵ�|�]ҭ���,;/(y�+��������,������(�N��6�6�_��ɏY�eNI{���ֹ�+�(��y"l*l�"W5���$�fy�s��[��m�}��xA�����x¼��唶l��k�׹?;���+T����N>5��%���)O�l��g;F��5�x�u����[݋F�ͺ�	�T
�D˲m��uu_�wn&�QG�˅Gu�\�q���b���M���j'1��܁�YK��ҩ��'a�^��^G3.����������r��������A���2���eWq3F�/j@�V�����!�Q�^�����9	XA���QO?�-����X��bZ���U-��r�?.��{�=]f�)���sn^��k۫EGr&���M��<6l�4��kW)3+���ڇ��4�r�6��b��}� �;lY�yݻ���<�^T��^TkVҝG9:!bVL�?��V�-��K��v�`�ԍ��ŉ7)��}6i�J�@>�]5��c4�ː5���tw%fx�JD ��0BXb�N����V�I5tka���'ğ��\C�RG��ϡ�G��0�����/�[b��K����	'��\�R�����������D�,q��l�7o<C�3:+�X����2=�`�-��Gu��|��Pvx��t��(���x�]������⧟¾�4�J��|2��Y�o���T�#��/cK�?qy�s{�mA~�i���q�i{�;I�t�ƀGAn���>nE�����仩�o?��xM14�R�*ȽI�K��|V?U:.��O��8��3?k�}9�X�r�ܡ��K�t�?[�h�U>�~�bp�i�Q܇z�rq���n_��:B�G�M� ��=�B�&�b��f��.����QCp�G�Rr����@UC`�䶖�k)�KwJ3&sa�X3�]_z�y/$��7m�R��2�jd�)h���Ae��(~q̐=�w���|����پ� 0���a!��I���O�,t�j��SQsHTO�����E����|#g��1|=��������?UԱF�6,�x��|V��5�oWď�+�N{C�O ��"""��3��G�vI,\zO<�\��~N����+6����_����N�R*Gm&ښTJxtp�0�����������ALej��4��\��N�Vo���鄚�r\��fC�--�~�ao!m�u�m���JK[��� ���q���iJ�,���?�3<`rtr@⣗�C~[ZZJ ��W�V����&�u卦8���!���Z��@~L�[�]�;b�s4���n��ė0b��������NU�_r�8�+1����Q��\�5��X�kUp2���"�m�{b>�V"������p4k�?t��B�P��+դ�Dt�4n��`���(�Л��Q*Ȧ��ײ�A	\��p�@�������W�<���w�4���ͽ֌Pb�G��������S@$����k�垺K�u��[}Ɲ�i�&�u�3?������'����(��
�z~BOAZK�[)�"J��[xL��I���s�,i ������������T�����<U�ҋ��Ї��V����dϐ*r��&4;;�junD����Ld8\�jPB���v�A�+���u"|hA��gE������7Aao1�>Z��!�+>����L�f/)K�=v�!�AJ��O���,�W�p�T����`SV�b�R
�_>l�f�{��'?5M� i�����_�Ik��+�B9:����3�1���<�$8\�������=X�ͯ�����P�-�m�W-�D�6��@�g�<���𖯺c����?G�,��?%���V�"{Ž6̺#rQ��yq����(S�Χpé_bO4g����*OlC"8c��Q���!�j��;��1E��*��\h���[5B����L
�{���e��а�I���˾�*j���(:O�7�,��I*�{*�R �d����͏r��R�nk�e����4����	��QX�=�E{U��7��j��.��'����@/ؙ�K�Լk�"E��Z��
�;�G"w0�}1�0h�:V:!�a���c�_�&����cep�8��՛���2kh�[]___�T�a�Q�N��bl� ���h���i�q�о�m�:1��d��k�����[/2ֿ�`\���+�A��A(�M~�
D��j������
.��O��e�����Ԋ.8w��睇�!Q`�g/���ppe�G6����F[��6������m�6�Q��Pg�:��o==T$s��ML��.g�½!�7�:�	�M+x訾'oUxk�N���I�".�/O'm	ǣ��m��=�
_�]Ѫ�{o1�+H�~�V�Yո�[��z�:8��
���:�-�}[���+M�s�ᣛ��i*G�˓�;��Z�%w�����Y�-3'��~8 ���J��0\��ڞ�E�&� �KNu�8b"�����ٻj����eK�"��yߑ��;4�{�w�?�v�����684�F�q�9�e_v(<&��>�B����IY̛!p5<,��,˳i�=�#��o|{4 ��ZAu�jbw��N��$�����^�����G�T��h{�1	���I�UXt���G3:�Zj�[[���ђQ�cM^_�QTZ���TT�����j룇&-ˎ����{��U�ؕ-;����m�d�7��W��F�.��UA��.��͑�� ��D\ϾƠ�[:5=���  �Α��`e��w� ��C�o?zI�P��M�r�[��D��˦�۳�$��8w���Y���n@_h�rXIԓ�έ;ƃ��w26c�Ėdܤ������Q�+��Ӫ���_�D���-o��>� ���t������&.��``?��-�h�Zb��s-CԀ$�X:\��P'�\����#�|����D��)��zz�SU���j� ��`��t��i_���LF����8�G����߯q�s�;r�^yNP�ӸR� ���q��z�����mm<c��,_�Q����c�F{����y_>(�s�<����l̎'j����TҸ���&#>�a�I���C��^��~����r:S����[ uL��~A`F��		�z��7���U�Ŧg��7K��PP�����f��H�q�j��I@m
{�1���ۍ1���X���&�q�϶�$1��j���L�
������J���Ι��by0B[n��&��>�,�E"�>�4ݙ�6GCwg�tXϲ
�)=xÙ �X�e�Vt�����1�Kךm@��:�xVv.ޛ�#����������D�v�W[6� ?pj�%�v6.��žVdzS^s{�8�𫨷)�ŀ��);����Vt{ښe��e�W��T_1�,�D�Iɳ]ץ<�}�z�����1;��¦�T^u�C���w����J(|_n;���B����F�n�j����đC<�>)���G�u�W&#�2qlT��:
�ꁷ��\ݦu �kB��ҋ���q���mQf'��ٔ�'�5`�/�3��Հ�1����kx>'�����5���;0v¹]|��<�/&U��}�۶��:���]�������0�A�������y]�_���,G�=����D���6�����d�A�55u��B���Ə�+����m>|�pitq��cؚ]���1���GH�y���ε5���<�=E-�;�|���\��yb&��N�����tS��:�ӡa^\ǫy���[�9@�#}7�¶')��:���1��&�\�}z(*&����Q��\ɾ���cd�s&I���\ӯ� ��w�����&1��^y��;Ys��v=ֈ�ҹJH���?������F}��]Ϟ=�c�%a�I��FvvN%x`����ҭ��1p>wSVO��{Uu=�u!�Սj���%������iP���_��bjZls�B��(.G0�.�zU-Yx����{"r����]�Vlv0VN��y4����d^D5V�8�&���hz��tѵ"�c�_��c��
<���\8�4�>��3b������%OU���kmi����.�?�r�d�&���@6V]gy���v��g��F�~��@����l���V"�)4��gt�qoHws�D�i�L{�TM���#:�ڼo�ρ��z	lJ�[_熽h��7SݩҗSE�Ӥ�wf����[��x~���v��9�P^�`}S�jZ�hD�i���JF�E�C^����٤�����h^����*K�q[e^+v��߷E�!V֋���߸?NW��f�G�W�7q��gg\�dK���9��W���v�u�^׆�~�2�^c���OW�M3�lM�m�(�
�P�V64��E|r8􊮘��!��E�΍_K)L���b	�Xn���f����?#U5�Q11�"iR&%r%��>�,�m�nF�ش=sI��y{P�������CR���{ͨߒ�1/���P������8�j�G�k.�� �2;�U8���;nw��z������'��1�aP�P���#����)�kn���$>��(�rk%�r�鋆(�>}��5וL�3wV���;{�/c`�֥����� A-�{�ޛ~���ٕ��	��8���������ɔ� �[�qq�������^�;�m@�K⧭xK	j7`��q�\w�r�q��)Ks�-�Z���a1ٝӜޤf;7i������\�M��ĩ̴�L����q9o���6�m�<i}��_pSS���b���Y��~�'e7=w���^)y�ߜT;��h���
R&�=�/�d���D���߁�%�g#����F�T�������V��k�m2D�%�fQ�_%���m:s]ù��K��)����zzzU[�?GG��#Nwu"�,G�{6�O�{�� T�j9|������y>�ϔO�&�!�o榇�7��E�(5 ��Yvw��@���I��;_58vb�]F^�l\F��2��Y���@��d[�{�'3��i�un���M׎�r(�֬�w2N�^U�=�n0ڦ&3-������1KGҟݹ�.��N��1���/�2c����=b�o�S.�|pa _U�����J���՛͵}��]S�g�|7ȏ��7���1�T�������m��ӯ_n^�����x����5����ޣ<~��7��칺ۿ�>��m��u�����ډ��7�1�d掫g<2`�KI.�U�y�z�T֫����`�?������;���ƪPBS���	.X���5��$��5G�fƭ,����@���0�i��h��T��ȕ�b�j���p{�2ngLy�1G q��	�^�P}�|f���J�:�j��qX������*R�Y�K	��r�[R�<>���"M��a�O\��Q/'/�R�����Kq'e�4>s ]D���-���3119�X�W��37��l�rX\⋀����ܞ�KߩJ�蕭4s&UHz�]AR"�/l�`ط������çR=.c�ymmm����i]c��M��珛�9��wq�=�p�%%�B��8�<��2O�� h��]�`.�<P^��,�ţ�W���H�ұϴ�l=�]�a{��S���sx!���IZ�7(����������#/CKf���K��-�k�~(��8{A�H|]Q>�:�RTCV���Xq�,O]511������̲�������.�Wn�	Q��v��G���h$�\F�h�=ijj�z`�|W]]=U�fz�>6���W�!\ⓣ�OAN���bf||jT79���-�C�d ������]7��Iu+����:�vX�"��>�B�����1�)�h�����|�ΝS@l��Ċ�G���i@�������mQ��Tju#��4x���P4�4�:�K=��0mV���u����M�z��?Hdk���l-�,��eKe1K��ҁ߫l�Z���� UD<�&lߍ`L��,u -Ҍq�Q����	�TaS��ȫJ��=�?�_�,��f�����a�dWkv�ڎ�A���ч t'n�9ȜR^i>z��(�Y!uԀ�n�$�`mr�J��gl����I�X��f �}��H¤|�p�����^\��g�K���!��k�/�\��L���Xb�_2 ���]ȨϽ�̴9���@}�w��M.133�;!6XX��C��Dk5L�!�ԯ3H.G.��l[2�/�2p5��D��U�VەURV.�,B���1����'O�e_����L���Z7ZG8��p[饐�����Z���t�lF���O/W��0S��v|!.S�1���E�!L�d��Ɏ�<Wh��kk�����w`;'���K�Ye`�?��D&f�e�	.��Q��@w�/1���,OE�W�JW�!�-g'O�<U?����;]f�K"��CH�uׅ��h}�=i��l����V��.�x�[8��۽��e�.�D������%��� ����}Z�-���2�4�B����|��j�`�Օߕ��g���>|h83�Q�2����ٰ��v���꧹��jr=��J0��R�l�������/--=���6y�|�JfVV����r����W�x��Ek!�����?EN>�ʞY�fe������}�V��d��7]�tؤ�G�N�ɠ�N�?���2�nI��ޣ>S�dd|=�pu�z�����5���}���O�uu�jjj:���,��vU��E�$����'������#�$�������x{jû|��o���f+�p��:���,5�����s�MA,"��w��_�}w�����d	�S��}�w.�=���l�H�Z&"�����d�~���}������%�:y�B���~0�y��(tL\�qZ^Y�x8"�E�!�~��,�(Y�o�cn:	u՗��Td�nmI,���57�����9{x���Q������EB����˟�����(8[�[��A�豱��|�)�� V�����AEN���,?���O ����=�8�&�4�ɞ~�:8���qΊ��cà��i��[���,xg.��x)n�����%�}ڵֵ<u�r�;�WJ��`��l�Z*��"�$�����3S�΂�#�F����̬ �־~\�JKf�k�w�����p��p=?Ԅ�#���O�Q�M)��h���#��"�=׈~�N�|������V��d�lg����*���ٿ�f�_�;�Lm���v���A<	�����uz(�M�W��$�T��o�o����#�55q{p�Ş�k���ZG�@%����!��,w� �
��� ��a]����H����)���T^{,2���������m6.����l���#�SZ�M��0?;������۽8�=i	��"ps;���g;:R�����!԰( �W緁�1��oTH����Q?�|V[�x�ؾ�C�;���CEM�GA���3G�>���CD���ڹ��ǚ��1�"�����U$���we0�+!�ّ��HnTG����O�\�u����]��;�����Ilf/���@T���_rAt*�d�X7u�8�P�1{�r"���҃|�+k��l��\���EMd1��C���������ײ�rt<:�TwZ��B΄�Uq�IڠL窈��(�t)�:/Z�j�pJ9��j��ׂ�¬������K��b5��VxE'#r����84�5���]�L��Q���4Il�p9󅊓Y��T9��w�����t�)�#m��;�;<&�L%|xH�����Cv&)I�mv�gjXa7]��1=��#�l�±o7� �sX��&M���C�ޑx��c��WY��5�ޏR�7m%id��
�!�_kVA�4׉��,��]�u�R�@{�I���x����8,lI~9z��^]qp�$�ͣ���78o�����d����g��Pj�
�K�D�}pg� ��X�"�lr�"_Ѣm�韴T#d��KA/fI�.�|6&Ue�r��%.�T�Ti s�C!���w��t�>�x� ^f��
XK����.'��ܢN��Ng����%��r��n��G����O�U�u��Ύ���e��|�JUg���gz�:����l@����ظx4�:�u��%yB�!.�R��J��T���
�%p�w���e  �i��(Պ�CS$������U�Wu(jn�oܨB�5����Г#�	+�k�������P��wo�(��)��d�jW�x�?�[�6���=cZ
!���F8}��H�=���TO�'$2�z���*����?�VA��@h�C���c@�{oRܝL�۲[�<L��[�譊��E �VL��Up͡� ���d�RS��*#�>@�o"8�t_��1���_�wxr{�@���GY-E�N`j9����N�|��_����Bk���A$t|�j���v���W"�2N��sﭏ��{l��|Drܛ7oznL6�~��:p݌�����A���^J=�;w����+*&�z��f܇���i�����QI�r=(�3�#}Mxؕ���$eh��(����fQ�,��%�ث.�Ш�,��=~�AW���B!�{Y��)k6_<Α��[�ML<�oʿ��ɓ<����	c��>k��m"�KLL�M9H�1��r��P��/X��?2��mq��_�/T0���������WS��i�Ke)_T�X�� o{�.�"�>�Uz�T�U��x��i������#|�N�<���w��{w���8���e�b��pA�.3[���h�����j�k�F14F	 �4;+�<�ya�cV|�%�$N�!Hq�լ>r1��#G�J@ȵﮡ�w��l"B%��^��W*��P�z1Dqt�>F�[����/pT�_���n]B^ N��1!�T	�1R5bbD~-�ލ��j���Ji�Ԟ���C��KX7��"��<�[$���XZ����z�����ݽ�x���vu}*����h,�u����+b���aϸH�i��A;�|R@AO����z��|��O.�ǀ���
��N���N*8�/�����ܔ��}�/�؏�y�n�E.[v�M:,�&���`k�m�k��K���T8�'W����62q�Բ���tB��]���^��>��I�(HT{i�aib����Kc'�Ͻ����j��c��i�<��A���ҷ���ڌ�_�``�_+̻�d.^�1n;� �m��q����TC�,�k&,"��u�������ǒ�`j�5L���[�$ p�^�,Q��
�b�{�F7:ÄVG�_�ɴe0����x���d.��]W�f�#�2��;���,�$.'����@g;�q-��cء��2yڕ���#KgR7�����&�)�%u/���(S�{Lv����l.��y"��T�o���8�x���MpPA29Q��M��>K�����'��u���O	�K@��
}�;~V.�*@>���G����u�'bY��zC��.϶"�(��+M���B{"w^��V�A���KR��)\�ŉ�w�s>��+�.�n|�nBE��'5ϸ�D���8d��a(��IC�|5@��:G���C��.�O䟬�	=1b�Z�0��' �B��s�wԧ�{�����"#����%���qe�q d_4���g��m ���׏��޲R	�)C1�1_��f���r:;;z����U��%>?��zL�bD��h���bMLLd[���3��;�P{���8��<}�����R� \��`���c2�:��?�4�"ʽ�Bt������u_�3���w��ܛ����xo�*��m�WI`�����ﾸ����W?��X�Y(Y���e@/��yo��S�����vޤ�� ���8�q2��-��=����t篡;ھ.G2��u�o�'�>qr.����k�	ۚ�e�ݵK�s�6yް����%�� }E��ؚ�se)Q��~Y��<ʟ/��/o����5^C?�����E��~sc\�=�dt���5��}-p[������(���]�d��A��<,���W}��xh��q�4��]�aF�y�<�|�"�́!�c?����1	�ac���MGfq$�7
D���-�,�W���jk_!Z�a��p��}�˓=;d��W3N�����9����v{Y!3ߢȸp(�:<��\�|�ߺ�"i�&?�zo����z�i3�WXޤ��U�:��-gj27	�s��
5N���ͺuX���ҲM��r-��
BRv��Vʉl,�6��&�����>�У+��̼?ނ&�`#>�؟���||���x�ΐK�U�6��ߨ���T��U�y�m����郘E�&b��3�����qi�e�������_�s�c�>5���>�x�G�i���|AҒ*ш�}�M���ܣ��YA�*�9z�h$��
6�QO��P�s�=xF;�)�ؽ��D�5�{��������P�ˠk��P�;RO��b��=��[���Y|@*+��?�AG��ׇ� '26b��S�znF������A��:MC�ȗ��2'���9���J�繋��1�.aKo�^;Gڋ���șF71ӑ&���'$���W���|�����h�7�coM(�p�[��H��W	=���i�g}�C��D�O�������v�'e���s�jTLw�ܴ�<+�G�E�1,�A^�=O�߂�^"�MV�?�7�&��.Ad \���/�$��Q�eD�s��&s�#8;�0!�V嗫b�e��p��Sz�ެ���)��L�ʋ���wz�=�T������U1�6w{y�]Z���d�n��D��g�r0{����?k�q��ۄW��Y~ N����О�Xu�n��i��	oIy��r�.����/�^<=~��+A�J�_�	�����{�G0�'����۴j\��3��6O�$����& ��Z�7p�,����1��2���9�Jq�7*[���� uѷ	s�R�|D����M�1O~t� ��<� M/�w�+�&=�!�ܽ�|5�7��J�a~�������\���<�p����m�,������fy�ٗ��$k�h���D�[����4��������$C<�UO����m@�u���u}t�<�e�����"�Z	7~xm/0S��c�@��&܍�B�<���%�.�p�?����"�A7�9��m�:ٹl����C���te�4hkA�����2�jw�����)�f�����ku����&�l0� d{�����se�wy(�����m6�v.��.��l3��v<FkN4==�>���� ��9셍���b��h�n��/���q--�|�r�D�â��z�D�q5�0c�d��/�<�K�*���ᴩ4�8�"���@XcA�<p�3C���0��3iqx�IsE�g�A�#�ר���(�i���S��������g���I�1��m��A�_�`�klJ�㦌K�l��70�Y�h1�X2���^ƬX]��=�5d$3j�0c���hӿ��ၽ=�"�C��C�h�h�	Ԭ:���嘣KKKe���g�O#l�.�����SR0 0��g�Я�l��LRg��(yˮcH����,F��i���Z�q��;d�b����<����n���s�ܡ&PP�8�F=��k��o��p2{��]�E]��	�����G7 (1��{i6���_:X�'��䙥�u/�#x`��z�߇o��W������~�;�Rjz|�ֲJR���((-YS�e� b�]�*��/�Ik�n��j8����^���14:Q룜�� ���Ǫ�N���������b,]�1,��#����yӊ5�}_���U���3�K��?S�j	���Ls:"�y�0 nk�E��܂��X�T� o���P�7��p�a�T�SN��N��=�>�Vf4|4a�����L���&��J�86��%�8�)�I���-���y���<��֤�i�0�Y��@��^����u���2��8�<��x��)�rD���e��.�`t���\�$ڏ��T[8�^������7�V3첽������ruNZ:����CM���[�[���cEi&h�"�wê����R�@��uh1�a���7��\p��묢�;&<����G[�W���9ý�u�����d|!]��i꺹r��YGiN��^.�������[,���|<�ɵ���e)��V>��u�v��_��W�GQ�3E���r�
���d9����m�N��n�z����z48v!�}Te�pB���D��=�z2{'P�*R0����B�.JݺAUa�3?�V��
������DP�[��^g��X:�ΰĢ�Mzu�/��ͳ�G߅Xb�V-�UC8Ƥ�#eoOSqkR�1˻��X�?������5���<4�l���v�4��b�'� tvnn��RȜ*�7;܇Q]��~� �b����䛰5;�
�����x~��l$t�T���$��5��坖uI���@'Q:����l�ʴv�_�ت�.0�f�j�@^�o�m�.$<}��%��y�Ȩi�T&!���-�J@սT�D���I
�FL�T7+��'�-ɽoU��F�樨G$ O))�=��~/$Z1hM`������D��P�����2����4���;p�[��{�g����A>1�=i��ۉ7�iFL9�C!���̞Yj�P�5e��L�F�������-���Pn�Nx�GL0���}��5L+mn����x|íb��;K�D2�Ġ�p������F_�Ah��'w_�����Z�T;�������,�8X�,�>p�iY���7n�i�/7??@�t�a*!�P!5�p�׼Bs��?��s�jNf�ϕ�� ��Ƈ�9��X�� L0�J�6�F�����rmu׉g~��"�7R(���nhDۑ/g���dH�@�)#H�;���k݉��_U(����n��'M]��a����]^��'_��R�M��#������]t}��aC�hzz c?
�_�wXH^�.�ዂ_�9��D.l�J@>�/�}ت�V�4L�U�=j3$��&T��,t�ѹ�o���[9֝.��/w�U;�v��s�b=8[�♜7��Q?V	��W�U�Y�ZP�x|��������������?��q�����>��Nc9q����sݜj����IU󳊆�D��	�]eQ6�,x��6fLc�j4�/i |>ln���D�aؒ�l�����J��1a�Tˀ�����Y�*Θ�ʾ��m�^Jhh���H�詈�d�j��O�����R��K��g"h���s;�i0}��u���>z�W�*�H�Ɲ'����h�s�o?����^��@*�%�E�{_��mddem}�&�o���4���YW_*�<iP�v�+���o�"Eg�)E���M����KY�=��?��R&�4"}d{�����7��V��c���(��K�������l2���d'g\* ���)mU�Z ~�����VA����;�Ʌ;3#��
�s��&�����\t� �q��Ș-PX�|���ѝ"��ՙ5�ض��ԟ��%N�뜞|� �u�x���D�d�����Go������	�������{�����5*bz8�eb���R"�0ziQu�����0�Q��b��H�͓�������.��k]u��ǝu�KW���]f~����Έa��tI�fq�'��/+����&����q�44�׳z' ��mUf����0W���!�z[
�H̙��.w��d\���#�>���JJO��xlO���Z\��cߞL𤐽{����W����f���(^ߚ�<��vH-/+���$��n���[�la{�o��{���%r�OY�?�v|�F�?I{�B�;~ ���[ѭ�q��&�4�o��YjF���g��S�r���Z�$��P�2�Շ8Xji��1IvĿ��67Q�t��ͻ6���͓D����V��ǭ;��E4�S.ww�i��?,�Xv�V�*0em���uu�'��}��*� E��!Y�N$X�#+:�=�F0D�K@r�I�Qr�#���pw|K@�Ge�����x�����(!��E�M�3D*#YWF��q�k${��ɾ�.�ȺHH��^��6���5��V����xxؗ�=�s��u��uYm��A�|jt����D~��ƛ����ƃ�\~�'�|JP5��6s�����7��Z�/ �d��]8���9!H����i�'����)ke���	N��y�_r�&�6�֭�mD��zд���=P���\�ᾱ���ǈ�P�ڥ'a��ͭ�`D�_�4#7g<�i��?`-��}a5��>�YO@7����<\���3lMm��`��S���*��IZ�6��8����W��ԉ�l?�	�^g�Ҫ�V�����H�ݙ��sÅZ𑉷1�S�
6���}<����O���R9����FJX;��L����bV��ٚ:�/xM�������M�|t"{���gb&S���te�Ѯ�P��������	B��,a%���<��)Hp@���~<���u�����NR$g���n :��4���bT햹�2�+5�'��~/�d��~��E��
ka�Z">�[����3z)��:ŪkgG�Q�-<�J^]ݽ0*��,��w�����q?b������}ݣ�[�nǾ݆i
j�J��+�%7ا�����Qv0�~~��+Z$j�p,����H�}�zs ���p��f�K����޽E���cF�{"���?�>�\�?C��5�X'�%Fl*���7>|�A�*��ھ�G���������O����Y�:N�i��;o�4�F;@IJ��򒪊	��s�
��	��z����y������״�e��h���f��FFc�N_���fV�~l�me'<���Q�qs�JE�༎x�[ )�1,����ZgbW;U^�1V�Q��H��8�S%�i*|�'�����eC�G�P�p�5�?��Tz��-:6L�UT�;	S�;�۱��)���=�D@�ږ�`���n�-����ȁ-8�:�܋u���~U{s�k�����NA����V'\�U�w�uL%�yLF+ϋg!"q���7�Ŀ�0E��U��uߴ�}��염���vOZ\@o���~�ư6����r9�HzT���k��9����D�I�N�34��-���8��N��NDT���HT9@��&�+ۋ�̧|���Z�H`ܓ�#���-���x
-�b��D�I`�6��{�B	�K����I�3�����^`)-8t����6(�E%�29y�OD������U5�~*RI�RG�	�w�6�$=�&2x�pKp�ޙ�24r8eLz��5�U3Myp�x���x�g�������F�B`�Sr��Iu=�fE�ӗ�I�'�����>���� ��9IK�g��y��6̜b<ot14xϘ��C�[ �Jbr[j`���S9�ן8\�aY�Nֿ�;j���[ ��=�\,�>kx'QtZ������|�;�u�
�R;~�Xo�[����K�"p��b8KMH<���)�K�����|����%���+�Gx.�&�����������zߑ�D�n��`0;���{э�?���F�TLY�_׈�v���>`y�W�������N��:3��/D�7U�_�n[b��zj�RA�g�F�����~���]�)�ϵ��*	l�da~an��7�hTy��^�g6����2xn˸
'im�����a'i���3g�e���`��͖U����$�((ɠ�r��S���U	.ٯA�b�6g����/8�9|���ǫ��n�%�7��9s;�u����V5cj�~��$��R�3B�V8���{�éhu������c�掤O�=��~��o]&�p�'�:H�{�ǡCM�IF?�0u�>]�����47�mG[ݎ��^k�>�UJ�������+ˋ�mǢ��z��q����oC�����v���jfEܽ�+�=���|�у��^��_#z��ܚl�Q��Ͽ���x
9^��� �^����V��gNI	w��ಌ�3�NDssW������2(k��� �i}���_�sC0r���y��� �d��~�5*���1i~�+u0������ s�ݴ=1��u]�z_�OD�s�Q0�y��n����ln��e܊�t���zI�#�~�$�k�g>�� t��ڂ�P9�J~�́Ć�h�2��lFcS������&��c[��.�G�Y��z⹀�Ŏ;�k ���o.�� �l�-�(��d�Q�y�ȕ���7Y�1;�:+&���k�"�V���z{�T�hJ��,{Ȓ�F��1i�,I��Z�~����0tmn��H�T�QϠ�2������e^�m}��V�B3�#�r�1$i�ۡ�=C,!Α���ځ��p���7���ƛT�S0�XS�����*} "���f1j����=@zA��p�P�������:�ܼ6����}VW�ɲR�S�u8r�7/f
���M�	Y�Z�B�ùT۸�C�~�%�Uܙ
���ݾV�v*�l\��G���?U_n����pV�]�LW��y�p�6�y�3��TGֳغ�������}V'�b�=������ ے^��vV���q���F�9\=]��Ǜ���:��*�m!턶u�m`\x�^�s�J��k
}Ѵ�Vɹ����>Ҹe>fW�t/��6`��^U77+�z�DMMmKH� Q���)�n��2m/_;�?��Ư�hٴ�zr���f���嚪��6fe�c	������c9}�O���d������	��P�1�B�U��Л9�Vg�����*  ��K�k�����BTTT_p�'�+�R���+~���+�>�Z���~�*..�/۱��m��-,�L�"��z
�D�5ɪ�h5 _q�+//?�����N�ş��̍gc,�认��CwQrq�q��Q���)�t[��)nf����f2���3^��m��UNp*|�^?��qb�CÛ5g��.���i�c��"~ Bt\��B�I�Ґ��V�_��u�֚j���Ό6�)�W��Ln%j�/%DEC�v��n�͐F���$�.����}sf\b����
3�9�[R���5A����$���GMVI�N���-+�B
�S8y'NNI��z�
<�p�����-���?�N��S9�v��uf�D�;lλ�o5�7�R=~5��
?gH-�8BM�qs�Ip�-����v��Ru�Q���cdB�A os��5]��ocI^7�Zgٞ��V�=��S��:����˛�Ξ�}��+����2$�#�gK�m�~��U��2�J��GU�0��:�����J]����M�2�<��؄�G)���Š��3ζ���BWשX���l�m�=�2=$�K��������@?�V?�m��~Rv�{'B'm�9؜i�!sn�@0U8p�dacc#�B�É*�����l̧	�}����������ߗX6�
�^�����1�R����#�W�9���`��Q��>�=#*��X�c>�x�����b+��E�+�<�:�<0���@;�ug�*��싞�����l�:\[��h�8�d��v�K7t�<\�A>��i6d��q��$]Ӻ�s������J*ԋ���ܹ��d�=]���.�jv,��%]sY����C������q��B�l	���sQ�K�9ʹ%.<u��������Qr��4)B�v��=���n+{��&��2��7m�L�m�3b�ʶń"�E������Sљ��AZZ����z�ӊ����DYTLlع��׌��羅������!c�Y��������jDsHp�:a|����8�������RX��y��́�'Y��Y#'�"?��͔��4�*��x��6݆�I���RYYy���8�tB�����M��v5rI�4��yi��7�_f,y_�/<}Qy�
շ��j�`�׈�/�{��s��9R&{�g]��t)�W&�ʎ
U<@tF�Z�o�4e�!�����nK ��e*_���8�(#���*N<_5S�����g��|����X����G���r��*!^n~O��/�iw���T�'���2�e�pu�fU8��7c�Z��S���=�O��!	��E�S~e �j�͎�OZ�w*���vǣY�=�Y��	Wם��f����IZ�1K�A۪���;�n���Dz���e��ñ[��c����Ӻ� ֺ���S���ӷs�(�3���*߾�da�]�m|�,U����CzfNM�hN���=$�8�{��rȵ��u?�s�z�����B�rӕ��H{�y�VPљ�洵�32�!FGS[  ��H9Q����	ݙ�i����g9��������@v�l�����J�v{�\f��k�.����,,���ݲK��6��8OЁJR�*����2���b;+ߥ���u���=G�Éҕ��m�����RY	��fj��G�~n�z�:��DY	�@g�T�b������[	㑟�nm�\�8|��ƙ��On�Vf��x�d�c�v�oL�b�J�S� )=n�R<e����.η����1�k�34:��m�;���S�vf������#+���e&)�E���ǲΩ[���0�z4���	|��^�_/=i^1�Xvd��c{=����|���l����腶S���ں�Ku�����N��>uW N]%c���7�6��/IS,�.'-��Â'�� �k��1pI�6UG����vO	
���J}�5��_w꽿�� �6/��;e�5�8��ƿ�K2��"��XU��e]8�:Q�xM��'����jZ�jh��j�&D��K���S���G�SAx+� �kڔ�����c8��õ� ��yk\+�[�(�3����N/g�7����%ܖ%c�Wm'�w)�%�g�Bv0����P)W2�nc��Ґ�]wrDFޓD��҃R�h,�C��g���:��O������i��B�,g�be�ј�ũ��6.3T���׉ �M�%�_����<��+��qJ��zR���y�'?�G���E9~��բ��U�cK����������Z)�=I�p*�EX��P�cojaV��M�*�#cD��&"2퍹?M��Vt�aʭ���4�o=����Խ<��C��&s�Ȣ�5�����j�p*����/�b����g�#Rq։���$o�����6���Z $O�S��:�hy_%%�� �~�B	���XP����Tu�v��V<����LIu�]�e�{k�����;��Z�	������1��R��|x���3_I�1���[j^����6����8�*���-���_�2t��[��z���o�@8g�ž��C�8�RܪSe��RK�r��M�S\���qK4��������MJ=�T�+v|�Mj=�b��~#����� ���Wn��hH�H�ib�B0�G>�ͩ�,1v�����b/���߹������J��/$��S��Ho#�7���ܵ��_(�e1P�c_z���+CZ�m�(SO!�lz�rЮ���d ����<����_�`J���N�0/O/}�T�Dv�h4�;z�>�a�"�\/H����jk�}I�w��Χ) ��v��{�6��4�Ѿ��Ѷ-&U�٭-q��tBv&\��b��Bi=�P��5x�[�F�	Ug�<o|z�b&�9��C�Y��G�q�n�|� 7���6]�El�סw�c�r�ǯ -�L��9q�;Y��۝�;<�}���6���Tn��f�M�)E��1�7
��tk6���:�Qɷ ���^�w�#�*����Wk��qK� C��9L�I�=齾��W��s��(~��ĩ���>�zrL�[V �e�㥒t�	N�gcN k���R�#��Eס\L�R���A�����fkv��\%��3>�8�KwbA�Q{���}���_n~~1�cRP�A$�.��Ս�RbЉ�:&�e�\�\�o�x�X��>���K�JH�!�}��Dj��+��������+�6ޝ�{g�s5&N��s�0cf(���hI��0�v�P��]!����I��U��N�vtU+*��P�R}�W9~7 ���XΤ9Tp=!���*Z�/���:����E��U��k3q������6^=�'Rʥ����iQ��<��f�V[�WZ�N���y<��p�:�u5��s��,wy!�f�Yb(H�!o��"͐]��r.q(W�M���5u��D�;�����ۻ���r.�n:Av/�ĺ�,Y�*-����I?9����m�J/�Gu��+VRm���=Hs�R����S���t�u��U�?��^�af��J�c{��:��8	TC{��C��u���#q�Y�'���g����E�~��_�SsM���C�iB�v��2�$�c	�����V�/<���`f��[��E�l�^�����d��H1�Q��aN��-F�X�hoE:�\�Zw��wc���6���'��ϧsm碃<��'�o�GM>J�>�#c�;�����c��DRH��/~����T.���%���M�v@�R�.O�Ӓ�`��cn����'M�S��ͧxm?f�F���/
�*�=�-ڂ��z�@ϩ$x�O������k��0_��z�����x8Ŝ���z;��R��� ��/;�@s��F^d�2;��:=���ykn�@.F�r �Sٚ����,mx�C7o���әtz�t9dc�%�3&�����)u��|����.�@����ka�#���^��s+�B�mc}�54�.��/7�r*�9܎�Y@��<	J����[7��pt���Euk�=6�:�%���������R��8OC#FP|���vqc�y�?!O�ڪ�@mԭm;#��*�E`��oOW����Rd\�./;�y>���zE��)�{<	�X�"-��n�"M��5�#�@��R5ᠩ�	�[X�&�3�Q�����H��"�Ӓ�I�j���M��~���%d� ����Y�(������ ��>��;Y@��lY���C���g�s{���Ar��H��c���Q�l4r
� �D$��}�]K�yʺI���m|��o��g�����S�������߁R�.��{�rP�]������~�y�������4�ב ��ڊ�l�4َQ�i��P�q�Mx��T��QJ�淇�zƱ��yV�
*W��'�Ķ�p�xy�mf�So��x[�l��������ކP�6�!�-�þ�P�AIP�� ���~�����!#M�џ�T�d�T�T��|�뎫��8%ů<��/��%�F̪�[��f����禔M�X�>�z5j����׍�v?[�����p��}Mp�U��F	��,S����m�Ej;�-G��n����������pD#����o�� |t��]X�D2޴]ІK�����O�4G΅�S���~�H�����+S�føĠ���:�緅d:�$�|�8���H���p"����3ox���%�<�s���Rc�ܞ�Q֯�boq�*�Og@��UM�F��i� ܪ��[��xe���	oW�W��s��x�EF�P���f�	�G�q� ���a�{��&�kc������=���XF��B�>�i�e��?�$?5�S���ތP՞���v��]dN�_l'�^p��c�=Z��\�+�;�6�'A b[Ĵ�,%��3e��+��&����)��؅Y� l���i�>�*#t�@>`�,�ʏs��s����֖�ɍ7^��١��z�F��~ϧ�M1G�!xY����G�D��RrZ0�p؝��KO�ޟ��h�
�.�*��@,ö1��Դs6;tW<@&,W��deeϑ�O�<���B���3\+���Ԟȁ���PQ�$ơ\�
1����"������������[�w� ��_��m6�:W~pW����� >���$�Q���$÷��ͳ���?�`�b�l�ܥ��3�Nnr�-�pt�옐����>��=
���J(�`�"ں�ܶ��v�^�_d*>����)H)���\�||�>?| ��%W��~t*����B�s��N�.��[$�Nﶟ��F{��B=�60�Q����[h�`n�AR=����@KN��	�o�5	���i�PF����S73���G	h����w�{?�zw�$;��������|^6��~g��O��b�o��NP3.$�>U~�i�ݵ@C_���j�
�,��7��y�pр�6���=�����s.4�N�_�]��2ͷF�I7�x��� ���2�M�vK��L$���u�Y��:`7l2��tMw�@�I��\2��}�+S~��N
���ag��y��r�*���tSs�����| �Z��լ��
$�8Ri����n�Cz�6�]�	��/Qg�+gH�mED ���!�5��Ԛ�LĤ5��
q���EJ���%^��	���m !��#����R.!{t�����5�[����j�@Y��K=c0^v�b_@^�_rmOY2�^��8M���g+kT�r���Dt4s$�6d��ں�T���:g��Rca�t7"��yxxL'_�(;���d>t�؞�!3�$�N����Ǟ�x>;�U��o�u`� ���)�L��ǜ>��D�u�W,X�SK7�Q��^6Z���q�j7�9=�)���� N��kϭ�ў2�@�qժ�I)�PSξd4�<���q<����������F?J��p6�PeM��v.3�D����Et�L�;�D-y��9���wd�)���@�+؟�T�{�|�u���[|+j`�oX�Qc��M�Ҙ!p�=����*ǻ	vN����1��?���G��n�neZ� a=�s�â��ׯ�Q."����&j�խ�VNʒq�t����r{���G���O��BE �[���4��k��T�j���௘O��
�;i�'�g�w)ֶ��k"�z+�}}�v�Tk��=������v(����� ���p���*z��z���K� RaB'�5�N��]�\�yr���S�?��$y&�4��v߂�d�Tn���S	�����c��7p�����7�ꅅ1����C��{xߤY-(S���d���O#��J,I���צ���|mƙ���$�Drܙ��������'r�b���t1s�k}�'���F�񌇋�68��
�������.�J7�xQ8����ܳ�F��1Vy�H�߯;z���w8h�Q&9M6�<�]�F����k,�-\��@�A����fk9� z_u"��a�wW��JH��)7Ag���V?I({�������{c]{�n 4�*�l5zZD������%A����Ĭ����Ҏx[@���$� ~I6_���V���d�������߼�ww�$�}:K��4-Ѐ�{s^K����L5��6gv��\(w||X$�}� � �z�OD��GN�я���j����{�#傋}C$T#
��\��aY���g�d�ͥ�)�1����NOt���4���lڻx��vi1�=��HEx������IԖ��؈��cf�70�Q<\hO9�ٻ�c�+�̳��6��N�Ɩ]��<���f!�1�"��/�aPcDo� �j.����e���D�\U���JD����E�\`yH9�L��KA?�NO��C˳��=�u7����ڻa�'��a���m�vª -_���C�\��p�l��}=��g���f���4K�����X2;&�Ű>��6�;�ձ��r�-���{�dP��v�b��SN����ꗟ���Y~�<��9"�0�\���>\���w��;[����S(��fw�r��Y<�,�PUJ~� dS��5�1��G��~|愞��>���o�io`8E�L��;�'�k~�w�=���D(q��K�6?B�׿�Zn��L֦����H�v�U���~���!��;��MB�����L�Н����_����IX�e��e�EuSk�W5�X�s$zt�J�Cl͊���4�e1�?�*���:�+����,�P�a��Y�؀���F���oT<�[�ne_s\���/�,��K�җ����Ir�i�}���^�����O �i�.(Oz�1!�g��>;�o�(-d�l�c����#�A�Q#�����ZO�*�	A�$R��]��l=��&)Ӄ?�4��2/}J���{� ����a��ۼ����i�%D��@�,�t��V#�(a����F�%Եf�)�l
�ߺ��@%{";���N  ��h����(\�
� X�]�ͯ��a�陰��&�!�2�D��x�k�9�5x�^<p�_�]c}f�<�P?�t��a�M���W���o�9�t>�-s��\ S�sw�~YD�	�g�B����)Zm�b�@�2&�X���)�i��w�P���<7�G��̚�۹����7S�k�ͯI
�@d�B���9V�Ց��q�e���2%1VY���c�M��1ͷǚ�7�v�c�+Y(�27�/�����!tA��o��l��짲����'�ާS�lz���X�g�(�=Q�;Q$%�w�e=�i��C��
3�jF�~��0VZm��.�)����ذ�5�ʮ$��,��V��0��JeX�"�u�!-�cV��M��:�����CgV,��ge>�<��i��ߠ=�BG���&��ty��f�xG����̐����I,X��㪛j������H��'��ǥ�>n (�0c(��f���9r�����7Dܖ]�$<-T�q�.D�rT
��opE�l)�(p���m���OW�޹��5��u�<��b��, �����G'ʏ����	:(��<�#�؅�<�	�:�?z�m�>�H���-{�E���e��t�ڟj6Dt�O�\<%�:�������{��������k˳��c�X�vln[`u�6&�Fb�HAI��Xl�ae��s�;����^�h��o������g
o��x��f���АJ�{�%�_����� �?�`ػ�$�[RI`k2֦M���`���gxO��
Z�ez迋����
)-��c���V� �_�g��rœt����hrU��3�pM��徘�~~�U!2*�Aj���H�7>|Si�|Ǹgc�0HI���!�}���OT���Ӳ�t��k:�t*��S�U��ƫr_į_ˮnr������F����n�r��Y�}/|�υtGM(]�?�[���R��SO<j(%b#,�@t!xR�-���Y��'!�7�	�����e���,'��A>yش���6Gb�&)�����{��7wí��[�-�tm����'��j��mU)��e�U�1߸.�"� K��C�z�[����s�'�l��;���}3�)�v�"��,:���Y-j��7@��k�����z�!| իL�KE����,�;�\ɵ@fD� t���VhS��=��i?}}r���:����Dc���%�'�Ye�s%)|K˵�y�iِ��	)'y`��V(Ab����
�"In6vp��,��eRe)�-�I}��'aJ�߿����?�!Ȳ��mS�'�'����~��ڕ"��)�u���yI��q�*fa#wC;e��w�V^NW�.�ɩ
Q;���
k��I'�W��
W���7��D�1��H�Ԍ-^�^l*�>d�*���{JU�@��ڒ����@0%$�İݣ7���ӭf6�����ί逪pt���8��:�-���՟��,�Kܳ�o�sJ{���x��5��GL��h�W*mF)�P r'>G�<�<b�3���v�(�5Ta8��;D�@��6�u�/$�Ig����|��e8�qh�i��Z�M�R4�ip� u�tak�;��Z�i��a�UwFk�&X�b7���I"�Eg�Dq��?}���C�a$�CfeS���v�ҽ��R��w4���������ml�Z�����[�A}�cɝG0����X���_)d������&�(��/�&I���u���<���^ڢ�{7���ZsA�l�]0%���h�8�s�P��X'�m�^�-����Wў�Ȇ͹�B-��A��1;6g��@��%l�d�׀z�@��fX�x��vl�K���,O"r'j�H�����<�~5��pl��S +ſ����w�V���4[ �fe�Ti�}tC1D9���)G������;�e��E�����l�{���L��Ћ��|��50��X�u��]I��K���b�\���_��
�7z��n��;�j,R�����<&C_OA[�I<��A��"MnC��0_�⤻�و�ޮAZ=��$%�N����19���ؓ	�ՋwW1�����UH�V�I��m��r\X_uI(��?����+)��*�d�壙�$!.zNذ����N=�ǫh�V��ϷR�������k@���!�jG��K* ���u�߾�$AX��K����f��ϔq�B/�p�ёE������WdK������	^`-8:���xl��K����*��ɔ'8�:!�������7�!_�v���v�'=���F���<w-;F�p.Et����[�����L-�%�''���7Ypv/�'VU6&���wR�!�)M�7��Y/��r��Z�V�\�_�~��?��q�?���(s�sn`|�$��6U�JX�z�H"7e�_�б��5�e��Ӛ�D��;	����]s���G���!�a�P�������f߂%�j|6�j�^p��%��R5�S�b����h9�j}����Ȑ����p��(g�Ō���̼�ю�g���E�ƶ���<�&͆���һq`4q�Mf��,yBt�a��+m�ڶ@�cў�i�iX�h�$�v�3G?���<A����e���'�Z�Z����F�ō��g��`f�s?
��]�� |�6��x�]��a�ҟ�����}���z����I=ˬ �չa��Y��D��*t'L�?>�棎���=I���	N_\~ݘ����v4�eSoHqDZ���y�z���PDU���5t{��>H�\*1����z�	�*"_�����L�!�����>��~��eô�pȦn\�֎)������,5�R����}�>��kI��kt�BV�ɫ9���1�;���@gvh@\�=��(��~��I���rOOʿ�����կ���߿��]�6����C��mY����������5�d&�X1ӄ�'����⥵����ݏϤ�[HNu��ѫu�!�����M�*���"�Fv&��������8><�/5�-l�[�m�x��c���!�g=0  (�*<��X�0`�(%�����(��r��w�xq����|�v�<o�J{�;�A:�/�ܧX�����Tf�1�����U-�� ɛ'ɋ4ck��q���������,�L���Uz�u�PVN�k�<���/+:D��ߦc�Ñ��Z��lO�4�`w++(�rzY@@ to��
Ao�<��%����>
إi�3WK�'�O`���I'���5�a�n��̥�I���7�ă���ݝM���i��+����SЩ�9��ϰS1֥�_����3Ks�*,��e��h�Kk�6'88�� �e�`���NVz�=f��������G����<���?u5�	���,,T�;�N���{U�R67�����6��A )�E��ޘ?�J$E�nZ?)C�e��8�&3�U��E
/��Kr��K��S�U�Kz3�Gi��o������&�/E8<=�b��:8O崹q�UW��`�o���}q�'ؙ+3�����M���ރ��߸ͭ��S�S���~��u.��.�R��k��H�)�륚��G��T��lݘn��[��<��l��+�*��3���=ϸ���g�O�GVH�6�9���C���`���?�p��x�rJh�|���S�h�aW~��.X�)4!���7���1�=�7��c�mG+xe�lڍ��伴gnE�K)�[��rV+�#x���T�\��'m��ڜ<ɕ���ѱ��X��Pӭ��Ŕ{9��H-+����5�m�ޖ��/}�Qqϒ9ޚU_���t̃WOZ���$C�g�_����ض�)�X+��(~� ʃ���)P�?r�$��_�$�|b}�-�Q� �nҀ��`[�nҚ5Β*�`sz6��`{w��{�e�|�(� 2Ra�V�^~0�3�xkM"|���g�,jH�`K�#��g�,�%�=���#���_�&>�A��O��RS&�N�1]�h�6]�zٱ��v�{��D�f1��ef���ᚚ��܂f�F8�>�6���cp ^p*��0jedݖɋ�y=~*��:E��'!#R��}�YҾK}�x}9W��,��'�S�q,�������wwvpڪj��.��~~�M+���*�V��J�����X����1�_�Jg��#�P�S�D"NPWBϸ{��&I9'}N�Z�_��DN�����=۹75�E��X�E	�ã��o��M��/	w+���Oz8��X��'nw_�,?T4����@ҳ��%^`��@���-������V�����#eecf}���l�9��t��T����x��	�Ϥty��$77��F�[����Ҷ�2����[�⇗:�~o6N���$.]ힱ�t��&� ��v�񙛝��M�!9���AU��Wh(�~U:`�)w?���A����K(�"����F�+�	;�9ztfV�k� ���֚9"}�	=NRH�����V'�C'���)�����r!��{\�d�t]��g�|Ɖ�,���sU��j|������M�)N�\S�hXKW$���C�(ljk=��u�I7vxl��@���qi�<��%�������2U"
���03�A*��'�r)y��n�yV$g�0��gF�&��)*vmo�4�(N�����D4�i6F�=��|)�ȷ=�̄��]nأ��T��y4�o������o��g������56LY��z�3��'��\>p�"e���������yR����u�H�ǲ�P�1�����`�Y���o�|X��I.�,�5��O����/s��P\0�F(��D��^dqdw�,&D�z�`��C��� �h���q��~m��hO�BS��C���]g����,�45$���jғ&/E��s<}^M|	^�l�RZ�5ڭ�;Bw�$��	�޿�(�X���iNi��,�D��TN�!��8�#p�]�Ǫ�'�J�.t�&��]� 4:ofB<@���rȪ�����ϖ���6��A�Ӭ��0��Y�#q#���K�����x�s���w��~cc���@�+ �N[�vͦ���.u�9�ۘ{Hm��xH���(��v!�I<��!�"ծyRS��
2Ƚ���.@+�䂍@�d_d�P��t��
�M��-���Hq��Sخ�5f��@�Z<ՏWK�+G:k�ع���f�^�%va�J���$��9�Wᣱc��J��
a�p�)��/H�M�΢��|���X�X R�����՞ڗ6���Z`�G`�%���� 﫥D�OF�þ��k�}C�Pg휳}���w�<��� �RϾB~���J�pF�lM�z��w�^���9y7�u�D~g�J$S�EH&;�z�K}�6p�k&UD��Kb[c,t�/�~6�
��3�_�w���<">��0�[}���x���N�E��b/�����$ih��O��>���ϖ�����u�ik�%��߬nm�8�������p��NL�݈ryY��p�	�`-��{��HQ�C���y@Cx@n<���<�	ߗ|�@:/�D>�M+��C7����#����qH��A�3���z�>�����SV�����_��M�|�gr�Y8�iD�f<��p���@�D��ט�\e������썴]UX��|d�-D�p%b"X����k��D�������Rɪ���t�N}�����u�������V�x��u�n]5�|Yp�VF�8�܏'L��F������i�<>>�}-3���<��&��歧kN�Jwױ�2f�GSC�xJ��� �K�
���|M�lT>r���]�>�S�ߊO�J����w\A2c"�`��	�R3R}���f���`��UY���+��("N�W)��?_�*��
VK��֤
�5��[��\R;u��%=�q����ɹ2]Պ�q�F?Deܻ���מ.��ollB���w��G-^>Eʰ�8����H��t��{s$^������v�*���r��F��o�E�6��b;���$sڷ�sD��cߟ�bV�	��~_[�?��;'���ˑ�?��#ۥH��i}�[�`!���g�B	;r�TsF����`/'dff�~�IN�o�C9�ݱ�l��[-W0�WhO9ŕ)��_%�zqmm��t�y�n�R+x���#-8��u�N�V���D>qS8U�˒0�2�ɥѵ��4�/��[�l���NIc��$d�V������im!UUݕ�N��m��7��^H�]8����[U&�k�`�3���I�Pơ�0-���L2�nVœ�b��Α�O#�
(�nƶ*7m�#�O .���8݅�(��ڎ�VJ���U	����`kF�؃;oi bV�ɘ��{��+p�z_���"f��fi��h��\����yQq:�/uU���p���.Q�D���LW��J����,��_��U��E|$*��
���&��v�� l_��݄�FI	���v	��m�gW�8�� 5�q)�B�����bDMG�S���e`��t���ڍA�|3���������G�y�|��\.w��*ɮ~N��w���R}��}��A�W���\^������@��*�η �a8�������m(�\�;�d�nǑ�vaF�R�n�O�Z����h�M&d7C����ɓ��~aa�YY�i��p:.�3�S�D
q���6P��s�K��S���_�E+�Z����`e�/�/����!�yQ5��5�T\�A�撩4*��>%zIY�SUJO�����������%%%�R��t����T�M����"s��O>G�������."�t#]���HJ����K����(JJ	K/�t
H��.%)�t/���������Ν��<�ܹ���m��+ݜ�U*��ӤU�4��>/!d7���,s=������N=����D��s���%C��͏��P�CS��F��$!pw��N芧r���[+��������Y�v����D��[9����\�A�dmmWe����>����|��s��y�'��<�tg�y���N]��;ő'A��#��њ	�� �N�w�(%���(���TJ^S�����m��$ţ�ǔ��U#i���+�<{cs��r� żK� ��@�C����#V��E��i�F_�|���h�vF�}f�m/��L�~���%����<_��ff��g��9oծ������(� ���2���D`�CP	UR�)����kǴ���f�<� .�K���(3$nB#4 ��?9Ҕ �Y�<3^X_YK͓>�"A
��9x��M+ �%'�Ɉ��=k���ѐ��8G�6��q���m(Y�o
�a�� ����62:�M��xՆ�t{hӝ<"~�g�m��%��fXy
q�X�����lz��O�?��!�x)7h+�u*c:6�����SuU�'�#���;R�o���A�G� ��?t��H��6H9��ʳ�Wҭna����<�?��7J(.�կ�o���J :5~��?�Imy�˹q���.*!�Q$�������U�"la�;����a�u����͆RI����}5933��'��X����zza�W��-#M~���60d����2a�ZfO��5��W�?eWQ�dP��~�Ϩ���;9 I���QOn�H�G���w��z3�=���)������u2���'hUm���v;�-ak�����ηtg��aDћ��Br���k)��̵Y+Ƽ��,f���<u�$�'�,g� ��_t�اII#�]�xj���]��ah�t��A�%W�I�,�4 e�rU�Ҳr҅�V{O (Y8x��YrETP�3��2���q-�,|���W�`}ǧOҽܸ^
��D�ԩ�O��)&2�D|�p���?m�����⽹P��ĽO�=�8jc�?�
}��ocE:ٹ���G�ăc��ui;�ރ�#�k���Ԩ>�Շ��d��&�#�v�ф���|S{3�0��_�i����qEk���8�7=�$�ɕ� ��~�lb��q���$���ؘ�bE�B�Gd$2A��t�vw��*B�æWUQ;=��QaeWi�r��f��*�-P�C�v ��ƾ���6+y�=�b�hSr�-��T_q�_��squ����Q/d���A���K:ܮ Gr�N�7���X���]�{����6v�� ���v:���0��+S7�J��1�ʻ>Z��FrK�*z�|��8����_'ߗ5�w�"kt�aMlC��O��d��mxi>L��&B��Њ��?Z��C��=�� v�߻ᡷ-�~y�f�X�:k.^Iى���sI�G]�n���XG)�Zz��'���;NN�aE�'���}@x�D����"9(��(qp� D����4E�|K���bW������|�0.k.�Y~��^B�H��~�<�¨|�(H���ɣ��7�/��Ytէ*s̟�O��xƺ��+=�`33�A�י��|��6w��!�H��d}X%bz�]ߠ)9+aO�&]�
Ĉ��+�%^�����r��gB��&S
?l���S<~���[�^�?�@�d�|TPƜ�����4| ��*�!�s좭&D�U�����e	f�w
ǥ΍h.��4ުCުH�}%�妡R'���^z���.��	�_�I����D�z#���r�E7�W���{�)�\ �����3��R#9Vq���d`��B��|@�d�����AP߿�v?���IU�7Ӣ�h+��������3�Sv�F(w��y�f
��eh�kF�;��{��J�,_ҹ����%� ��&hfN)9������2E紧�*�ԃ��KJ����������HK���E9���O+�:i�wF	,M��$@P�f u�L��Z
;s����7�(�d�Y��y��a+�4�b����_��	P�a��~maى���Uf�=RaQK����U;GY�d����w��uH@ǉ�v�]��CY�T��-��4|�K�x��^1���۵�=�����WM�$��.M'(��I�U�����yyv�@��=�<M/�aPnq}�3�����Ig�}��ϟ�6���ĵ��{����;��J�����	��q,Z���+
3���h��i�ӺP�=��gl�*i��8x8Ƕ �����z&����H���Ŷ��b��TBDz��a�L����Ǚ
���k��x>�\�z.<������F[�,��Ǝ������b�YCw�V���c�������t��jE:�L�y�\U�?*r
x$Ɵz:%1c��:g?��>����=-�'���$tD��E��I�GO�$<��� �����p�2�"�Pܶ�X����p��/��m�_�����{�a2����Ј��?i��,�P���]�^`���ͫkj��-l%YDBL�k�YN����O���Ɏ����:dV�1��'C�#嘉M*�:�xc�Fۘ���04�2�"�M�iRۗ��'�]��|\ҟ�di�7�Ѹ��jt)�O���̢K�A��5�0��qҰ�Sp~k���/�<q���?���"bg���u�P�yWq��s!������o=&;�]`��J UB���^�O 6����Ğ���Eu����}����U��|������L+MM�i������ע�F��̃�[g���ʗ=�ҘWnKz@����s�RvK崽�'=�h�h7�~��������������qE`V���+�O!AS����A��q�".�����_r��<=�c0drSS��\T�F}'�-4�2�n�;�S�$��N7__Q�l�{����>���˦��*��]H����|�z��L�~Dr��X��̚8PB#�ý�s�A���0�|��+D� �L�3A�5���g��5�}aa�k� ����,/N���NY��J��+)V��6�!�;^��7�L�pXe��E�ǲtX��q�t|o�~�jH�V��"S���M�#R�C������v�V_����!�5���i"�$�瑀ω�1~�l��U�~�qC����B��x?%��٤	4�z����+׻/V�W.�S����g��{k�@J��ʠdg���ɐ��J;��pq�����|���m�т>@zk��e.ψrB˳ ��^V��	��� w�5yrR^(���	�����.���q,��������zl�̽�TE*47�|q��N|Ez��y����m)��e�k�X����R�>�91
�i[���ߜHqw0,�֧�|:����ߟ�<���B]���7�jb��S�I��-���R�8�k%O�;�6�=*�$y,IIh�4
� 8�*��K��r:3��(y��(�LF�F�����S����f�`�_�f�6�]���0�(��0(�??���a6�28��b}1��"��c�X�"�Ƣ9�x����V����n1]f��ͅ�Q1���7U��9�?�f]I��!^�E��^���D��e �����\�2^���	�	~@T��.�4��v�3I0Q�7�ka����0n�����9y��������q�ύr�B���+�Y仓�(F>+����zXbzdjj�	��L�*	����!X�G�/# w�K嗦H�����=@������:׿�V��l3T�e&��8J��:M����]}�I�Q�ۚ.Rbv�P�"_a��[z�lk	�i��|�$�%�R�{����[���Ӌ0�N�v�0�Q+�U#��l�*66v�ތ�V��fo��o'�]@���W9�K�R�����T��hN����>͡���U�w:��2�S���2�� =���Gl����R8�Ks�9����a��EQ��'�z��nP�7���]����+���e��~J����~��	+��@X*���b��̌j�#P��[��)rξY��L�˒py{�C����U�i)����5LZ�ꬋ��`^����M�=C�����ќS����2�/p�,�]�8��s>���i�k �2c�@R�oR��#s�����U�E�S�{�o�]�1c���
H�_��+�<��/�v�N#A��a�	��'���Rv��1�A��'�޺���]N�ԙ��U�t]|��� �NL�Tץ����������{�LE�j~��`F��7WL�	:Ó�X$����"[ת�k%)4�P���P9T���@��a4��OV��vi�Lu|;����t �?��պ��*c�d����~��܈���i= ����0A8�{�+ŻK���baqr0SA	�E�>O�?�:����%���o��_��) ��97U�D�T��!�������S.����W!�,,AA-���a��ʡ���-�s�����L�y�~	����5jS
��N�od��kMh�</�I��*Kj�Fk(�=�׫_2s~�|$�'��!�euZ����D@�=���;�� ?v���~Dnf���i9cy[ Y��239r�f�zv/��[�1��݁_�E��e��8
�
��K�7� �ER%q�"��}���Jo�nE�*�n����P���o$[�/�s�붖Fz��5�҂���r%kٔ���^U���h��v�$���{�/8��yl����KD��E&x�0c�بa���T64��W�P����8�L���A�ǫ����O!c6�O8 =���KO�Q�~��VwT��kw�;�m��	�N0c�z�Q>3E�p=@�u�#�f�}[ΰ������I�N���c@�)i%9��rty^�4��K@���V)��cwW��~��+ϻ��~�кO`��i����c�Ba5�O�"�����z绋��N���6B����jT�fNg8�W��[�k�A�W�߃C��8��"���c�l��F7{�X��I(�3�x����]Z���Y�Ã;L��2�@P
�5;�HM<�����x7�;y�9�c)��j�
�X?WQ86t.��\�~�~ �e Iw�P/zIpx�w�D������2������ȼZ3�#�+Dj�-���Q�D���ŭ�`_8�ց�%w_��'�>�`I���""Z��YP�e��췾'�=�ߣ�{�����07�yF�K�9������	E�Ng�Ӻ���^R���B�tk����7���Ӗ?5�7b<6�!���)Х��fu-gV���!�3�1�}�D9��PX�V'C&4@�O�V�D=
�r���a�S�a�X�V�$�ٜ��|�Za&�MJ��잼�~�?��M�\�~V��''i6�ٍ֭��Z�4���D����I�
�K�S0�S�S�%��Yxy�V�"+5�����&�I׻��쾂LjOAb})�y��q��>��C�Ahs_ޤR���}'�u��t�n�����@�7~$_��G��NF%��;�T}3_AW=�6��OW�L����z����R��}[����P��G}��'�޳W�y\s:��I�IO;7��4}'��᳾�7|�W؆�VR�e{1��Jw&�9W@#C���H��G� ����tjJ����c�֔��Ov�p���fn����T�=9����Z��R�`\/��y\�wH}�j?���U�N��%�@�y)���C6����w�T�\#+J�m�ɽ�K
4�������
�N��~�b'�ؿ3��M:� k=�Fퟔ2�[��J8�U`��k��o[]����Qv�z��vmhh��z��_�)Qh�: �����!IlL����߇�o��J��_1L8
��J��ޫL�̣�p�bX�s|a��Tq��AՎ���{��l,���ߧ��zi�W��''�PC���C����
ܭ��x!���o��s׳���?H�7{p;KCތ�RU�iKL�N�yw&!3h�d��%^MC� �?{#�֣L�y��t\����I�ҵ4�>�pQH���H���9�|�N� u�V#��Z�R~pdW�l���E'���������?�����F�=���hV-��I�X{�Ի�67��D�b�cV�\3&�+��~����>�ݙm-��q�]����a�I��x�576R����]~�/����CH��x2�~3 �	
��rv�e��|#U~���,��H��r|�>�@�#������++*,n�TG1��n�77�������
�ٖP\\�u��HK�,����Z'346�K��{P�T�C�N��;/.���3��Z׊���s�-�M�훭��r� �!�rd�0�ef��I\��]pӒ�b �n��#ŒGY���fN3S䍶�|��\�[{���c����
�~=O�������+N>��\,xdu��Z�Q�R��4���~��� �O9H6�+��?['i�3��Q"&Ǥ���z3H�cI	/�����3,�B�E��FH���tI�޶d���,A3S��.�T�/�e���x���UQ�ˉ�ç����ퟥ�9�~O�� �PYWgW������G���K�����o�������nN��}�1���Yh0�z�5�r^"x�9xy)�U:��S�uo!��S���C 姫'N�6N����Y��@uuV:�uR~(������X�����H&Y�_U�����o��"I�S��u�������4>�U�4ޔOv�N����9��1��[__oPs�tJ����m�t5(8�X$�g��9&>9'��K�!d^/��2��05��xX.���s9[������9��z����W�K��qo��c?��=���N8�������`�\ӁM�����rv���]���U�{ɪ���eѩ�0�A���E݌ȣ3�!�s��5o�W��-�P�^�1ˆW��� �wSk��h �h33���,my)�jSUE�cnBf�%aJϺX�����?>[�-6��y�j��q�$%5u���up��"��
d2��u*��1\�,��I��v�X���4�N���J��L��,L\:���t�O��m��-�_����,	;���R��F�u����kà(���iW��v���]����5܂Q�{;54�8\O��fw� \�U���듛��K���e�����_�������egd���p��*���,��I~_��y���ȸx�B�_`���}|0�0�l�F���<t� _�� ߢ��ak���!��n��u���S�g����LO��]W<ovM�H���W���x)gn�U]]m��Է��i�e�\�>�A��F��O��=�h�?Z-8|�}Ju����Vl.���V�C����.w1���5�>�;LF~�)i�_F�sٛ�3=}�r_:Y�Ԇ���who�>0���\Lpq��y��q��{�b	6�7� ]9���q���	*�~���+!�ĻS�j�Rm��ǘ�"��Y�D��r_�+P��X޸�?0_avј 4�0��������wB�>�݋���ܤ�̵����R�w%�픈�봪pH�;P"J����k~�Yq�M�f�h���"�i�JM�V�e$Hօ5Id��#@�]Igu�)@�n$:Z����㐬0ˁ��Q]�̂����U~��-َ�$J떿.VVO��7�1<j0��~�����-��Vr6�!�a�S��i/�~�5c�4f�/al,���"��⽼�	���j:�j�kT3���M�Mr*��<؊}f1��<$�U�~���jໍ��+s��8b��aW�E�V�6�6��u�R�=?2�x��M����C
�Emu�ѧ_���=%��3.ӯl�Y�l��B��4�ÄOH�Ŭ�u��[Qxs�*�XF�����I,<������,7ifO��T1�=N��F\�s�Ie��-,�����^�qz�	��䋪oP`��OSÑ�3�F�����&�dP��](KF�(���m�cg`ȹd8�v|�`:�7������q���^n�D���@rK!��>�8Y�ڥ8���7��q6r���Z��w9�������z~D"�h^ب�uʎ��ˍ�F}�_T���%3W5��>�q�Lv��
��7� �����ͺ�(��،���#QO)�!_��Fo��/ˮpN���z�Y�F��9d�_�����ir5�"�L*�}�!����bɨq�*WV�s���?0�]�N>2� s
�2�S�6�mM]��ߚ�:3s�'��	lD��S&v����Zf�P=���1�ۡ0�+u�ό�����r�;�˙t�ΣA�3#^Ϗ��OF����
����~
�N���I��D���`�?��	&p�H~	���}A���q�[�b��:y�.U�6���'
x���ׅ�~,��2+�h�@����XV�
�����y�% (}wqʁ����,IU�QH&��UDЯ��웤��Mp����(��X���o��(]]wث����⫊��(�R���G��>��a���i
��b�����o��2�Scs3��%>���<FBL�$�}�<6�ۛ)�����_+�$��h�JL�+mD5���w?Cw�lW.�F4mL}Q�?�~�8�>E9�G��6���(	9?cH|>��M�v�@�MAِSKuI��މ���c� A�T6��	���<weSv�/���Փ'�� �^��4��mZ��5#-�h�tP�-��o�ow`����ԄW�ⷢ߮z�W[��tX��$����vǫV��MLlz���n�F���V���R������Jl���h�d���[v�/u��o�i�]zV��K�@�̄	H�~�NX#cEA�ew~ff��kYk_`q��R�/�|�-<,��/P�EAi�Sp/�7uE�50�T9��M/�M5j!��R����bfH�Qc��pH��i(7e�!�� &S��˨hu��:B�qH[�0M�BYO��R��m�ST1�ԯ��HI�޸�ΐ+A'��O��	J\)�����`:���a�H�Ϋ���{�v���1'����s��a�8/nK,�{=/@��`�4f!����c��M�Y�"D�n�<vs�?8�?Ľ��� X�DM3�مE�39ʒA�_�vM���AU)_j�OX� nIE?�*'���������)ۈ�����y�ۍ��Fl��0-)z�cM��?�L����6q~A	K���W$'�A��T�լ;a6�N�s�[tV����xL���4��E�!��Sl<1��gݨ3��k���а��03z�q�D�̅��7��ք8}0�&:\�Y�eF,S:~������x&QrV7�.��zq�����ܬ(�eA>�"��#͐>�T#�i�HB5u#4�,�n�V�u�6�:�����/p���z�t!4#rG_����!�ɂ�~��z-�u��"� ~�a���r�/�Y�؀p�WElU:K��NھbR R�C,M���6`���<ڝ���j4D9�xjM���y��t�8�+!�l�m��5?�[�|�K��:�}����vzJ�����"fØ�F
��ϽI~ҳ)���y��b���3��0{�Y�WލT%�^�~%���m�����3{��H?�½� M�uN�!<Is�#7��JE! �(1�#奓@|�UݏN���k�'!�]�c�_��DQ<��<S[�|���d��Ӆz�j��J�C��$3Q��r�=���}�w_�EQ�}Ѡa��#��ݯ%//I0{�oH�����q
�v�:�?�t�"`����
௼��F�c9O���/���܃v0�h��x� ���j�]y34 �ϥ�α{	\V���SH�;!>#�,�N�|f�`Ԇ���8���^Պ��/�Y h�v��j+_T@��W)�
GuاoiL�?VCRA����G8x5�ix���M5��l���sNz���
~����>WN�-s.*f\vK���Ɠ�u���%%���b`+�o�- ��]HS�`d~��W����T���D��)el�h�gz��׽癛�?4�M:z{f����4�F���	}}�'�06��v�|��ڍ���z�N���F��^��*�a�mt&�S<�V 12��<�S�/�
}`��AF�8�35=@��b��P�H���
��O�dh"9A� ��hz���^�pE�#=P7I�٭�Yn9g��E	M�7�D���?��4��V-\�}�dH���_�=�
��l/A��|1�/����Î�i&P'�/�t�^��]:fw��^~�b:;���k����9�k�/�� �����^0tZ^����� "�#��i{�[��;���]J6J��O�(E�E���L�͏��Z5}���R�
Oo����l��p���i[y���I�c`�;��Q=$ƥN����ԛBPqbCK温�ow�H=@�zn�ޮ֨#�hs��@jx&IB&=�3�a�����}�X�*��ԭ�QRRo��C�t0���~�l%D���!9f�9�Z�3��a��w��2�nÈs?��)sw�:;-�Ћʉ�����y��v-��O����^����Qra��hhX��׳)���=r2��3V9�~��Ǟk�& �u!N���פ����I�MB��Lx�Wg����Y^��m�z|=G����n���(*��x����M 5��k��� _N�
���u���A��!PX��q� [���b�'٣��a��T9s��׍��9no:H��c'Γ�RFْ�l�����}���Ix��,������%a��ӯ�E;�hZ"���r��8ā`�I�tjv�����mI��
㲷>9�^V�]��SoY�.b.��Yj���l��>p0�>󇉀�)2���(��ӻ���^k�鱃Mj���d��� ���2���?�Ӷ�����Vr�{�C���;q�����g�9�;�_#�g�+KR�[�W�?�Y�����6"�$�Bd�Z�*�Ӭ~��@mo
��؄�֊��X���b���_����Y`B<�ă��FW�j����ꄸ1�)��̸kޱ��V��������h�}b�i,�5<O`�t{���ʐ당|�ԉ���)�i�\Y�Y�����]y����{���(�&�S��9���va��ڝ��x��	KKr���2�=�K�>�v���2T'��� 4G���T?�F��)�zq�M���VE��$�e�
F�_e�rUmi>��~o�pѩ2�$���A-�qߔ]Y)`a�/��L��'>��K�E��Ta�O��P��E!�2��'"y!@���L_��'���y(���'}����;9����؟�/;=���͵�e������8�B�`t�R
�wM�Z?[�U�v��W(�����F�W����@i��!��ay�[�����0=W��q�e\J���d�ȸ�a���WAo�q���G{g��R\c[�M^�>��@o�<�I<1^�`�ɺE:��n�����H�+��cE��֌w�ý��-Wq����V���{%3o�_�P+ao�����ݴQ1?r5$vss}~6�I������bo�z�G����q���_șJWJ�3����ย�GDj��BmS���+@�Q9l�KQ/"ԍ�.�ՙU8���b�5D� ^�"��w�1,���[{5��?VkC�n�Ţ�#��O���7������F�C���}U�҂�E1QM̽ny���C�l���O���%]�8�|��JW�ٹp��E�7������=���.^���my��=N��UQ�B�lTߖ��KcR�Xw�p1ԣ�A��.Ja����pzo#��i�&K��`d ���媟l�gGϭz`F��-�vwZ��b�_�'��k���5��'�fsw�2
�`-�w@��e�ט�$� ��͇��ݷ*J�Q4��l/܀�5ݛ�U�>�����z���t�������(��?�u�;"e	��qj���7(vS)�.��ʶ��:u�9�A%5S�P�bQo���ׁ������D`I�EupK�6���2���4�Jg[�l���*�Q�$������Z�ZiB*�r�91�iq7b�u0<�<�f2u�"uڱ�G;c0J�)hv�MGǙ�x(u�k�o�"mo�b{���n�!��L�gV�]��{A����(�~��p�K�}����S'�*B��4l���>G��.Ԇ�˷�k�E�t���m?m���E5?�S�e��S�[��_]	}y}�e_�jPgG�;����ț9�e]�N�3�'XI��@��Z��(U��Z37���SP6�DJ�8�\V��"=�$!D�CNL0.k��cO��툐?X�ϬCsJ�a���/#�E��݄l�l��vq��򉱘-zl;�LŪM�M�6׻��J�ڂ#��7��>�	V�p��-u��.�J O;p��k����ٛfx-�2o`s���n ^��ڹZ�ǯӀ�^eҕc��73����ڷ�J��r��2ɟ�|�J��?˙�Dg%��KWא���f��dG��3w:��*j,��r2i�E����]P�m�L���$�)KP&f���
@F�^��6CR���L�b�u��l�&|ѱ�V�� x{
"9D^��fG"d=�?�"w�a�&�G�%����Z��.]��mp���O^��=��Q �8��<�uN�؀}�2 l�+f#�m�:�ރ����J��3�2?IY��M�
���ne�/e�!˾ŝ�.84@aw� ������PVM����kO��^�/<d�N�5s�9N����e��O4�Dʹ���C�&�[y�D�@�[�(U3d�	)- ���wgb�A"����Л�o%�����>"������C5��]�N��b���ŇL����:(r�����%+j�,����SH-��_q�g����G�����m\�ƒ�H�tV:�5E���CP��X��c}��ƺQ�UyiA��an�ū#��+��R����u]* �{�: ��3cv2����bTء/�&�<�"�/eP#é	��+��UM2 �a�&�5�vb@�p�]�dB��MZ�)P��������2(��8���'E���T!['���f�ɪ'@I�X8`�{���@�t��A���[ǣ���o�9�	���f����X5�9�/f,/����]����f�J��Q|c ~��۰#< 6�pF�ӂۡ�I&r���ȇo�zxx�DL�Ɓ����*n�@�d/� (��5$��q�b��S����̤s�#�䝁�,��u�K��MB���-g����r�M���6�ۓM�p����7�S�hܦ��i�����g�1iN�fH���~�/�����LlaQ��L�.b n��B��i�UZ�0�i�_��~�V$�q��H]������EIxD\VXԣ����OJ���ǃu���dE"|�?wށ��[ZϢoR�����ֳs�i�7t7�	�-o48%�u����n�YH"�k�Gks7�6�~�)�� �jR���/�FP��ԓ�,��I���c��csĩߎ,}lo�yys�4s����4z��\tw��l>��6���+s{����$����A���!��ɱ���ܤ���9��zUX3�q�.�����_���n����o���2��S�Z-�L��,�%w�:+���O��S��BXi�;�����d2�P���t��X�R4��L�Q�/dL*�.[+�د׉k����n���g��&\ ��Z��-f,Mcv*��u9�l,ǩ"a �x���,��o���Lihii�|}�
�T�C��+U��RC�6d[���\GK� ����1+�f,wsiqY�[����	& �+l�
<�"-��9.b[m��[\��^m��lP�5v�$��;��'������U���M�����	-gK�W?U}�7��Z����BSO�Oa~�^���_�%�W
�[/���w
@���A�;l������>����6�y���S2�Ѽ5�Uv���ԓV���bh]7.Э3Ίy�?7�'��c��O��K:L�7;���,���� ( G��bo<����u~Ŀ�;����Ŋq{e�͙Ok~��avO�BK��yuKy���IɎu�s���A��Ϫ�G(��vC�f��#��a��L�^'�\p]	q�yk�����rצ��W=��s$W�jM�Rsӆ/��q�W����_�g���Gm��Ϗ�Zm�r3Œ�O�g������@���E�e� ����C�T5AT�"��@j�;�rx�qY� [�L��P��+00��u޷���-YdksKNj����,Utu_�>q|� 6��;Ώ�B��|yjFo+��*PR��o���82Nca�%���sF_�G:��#����rc,^��v��r���Q`�s�������]Di�����l��YV^A�#�����[�_-k1�@�{3��������(���;�ަ:}G���A���<ۅ*�N���~�D�+P�1@��o!�o�P�S�!��f��ld`R����ϛc�wv��]�5j����=�����E>r��b�&t֏�9i�[�>3_EQ�7_��46��ޫ��I\��F�Uߜe/����A��7���k�V�����S�Q��DkCC+���9�֫���`��������:����	����� ��5�����ǷA'�}�^�|{6��=�8D����d�,�ۣ��.::�����ͧf��c��v|糭�s�Yǝ��2�jtB�l���1Qr@s�]��'��焪�VA�ˤ��*N��A�r����hu�q�­s���EG6fj�꓏=c���n^CP�8��sٔS�����Y�;or?@k���@eOA��e}�'A��o���	���?����A��M���Q���-�2�m1]�n��Q���w�Z|u������͑�H;K��_��{�-8�J���Л��sް��wD)�!��'yo��Zi���
T�}�&����K2��.�܇����p���эq���������a�K�)un=5�Q}Ae�}p(�)ߘ�zĸ�Ɲ���UY�Y��T�5�C������8k��ě,�B	W_����=�����1^�~�U?�(�c{���7�:�L-~TGw��R��u���I����+#��d�T c6wa�e� A!vD���{@3����At�����ʟ����~�ũ�=ٓ!oU�ۛ�>�@�A��^��~���)u���O[N�8>@�6F��҃jbﵲ�������X����'�N>�X�����0�c���,���wCtV9��7��4j�v �_|Y}-tn����n*������v큸����V1a����G>v}�2bZ�G}�?˿����Ϯ�������0�N+�&Ű��҉*t}V���~�O3�Ker�����'@|=��V�矞��kL={O�Gh��%SdT׵�N>�yB	�0�`�v�����m�T��8�DԚm����S�_887���MU����F�o��!q���Zn�aN�e�@w8��[ҿ�����Y����R¨���vBo�%���yW D�!� �eQ*	�gi�Y��9���l��T��I�>O��EA��)��U����^��7�C����#[ǘ�Ҕ��{e��,`��rL�����t���Y�!"+�ɱ�� ���ڹMQL�B�k^�߁����5)T@`��n�8�'�7hZ�&�J��l����Lwd����r�H�{E⢽7���.�&s��K�;��폤A��=M�� r��H���Jhe^:���s}�A���J��e>M�I��E�P�^��gs���O���qv�`ߝ{��8�^5��z�@�D����nM��R�����z9��^�8�;�+��NǶ�)�2 ��5{Sk��9Tv��sӶ�=��[�B������nW�$��;�x��=�#8�Ы}����@�|�v7AVs̮W���C)�}�ؠ�����#���n����4r��$$�இ���?�k�R���A0/4Ͳ4�6E:� 9�p�fS����_z[母�&�;���R>>�ݱ�'�'j���6�E2���,o���H�Ɵ�O~;F\�_8��3|�8���^�`����ǽ����P�K#6'�r�7����a��а����o(���Rvo�w�02���Ĕ�2}7m�2����i�1b�qT�N�EO��{�gS9_���N�BdM~D�c�E��9��O�F���@|8X��>`j��k��jP�����+���a4n i& �4&�rs�z޳��̱\մ��>�ϱw�������wCYC%�����B��5�-�k�n���0T�ԥ��v ��}���I�߽���NR�M�k
�g�����:���t�X� E���^7'�r�L�f���8�{��wH�Y�q�P��mw߸�C��z[�ȿ�x���/%�Ma�CP���m`T���ז��1�O�A��/!������ 2���q����ivM�t~-%���#���i+�T���\ӿ{�a��kx��lnݐ�c�Q��n��q��ފ�_��b�,�L@B�F<8("�x��P��|,��}���ا���������`�M�IY��,��DN�X��4��E��.����*6sA�x�n�w�B��^��t���	�鬡ʲr�l��C^��*����ܜs;���l|@>���W7b�.�,l.����ZB5�p�z3x�ov���V�jZ��\�Z�<���ޖ�`�O�3�f��A���ֆ�f/�9��j��4��hNLv�$},���-����=��ٜ��k�Ǣ���L�tu�b��ih��ʷ��_���.Ao�%�*[�"Pe�+H��rߺ����U}�!�PO����Z�sV=���q���z��T*�L�Hk�%��hV����~g�.�����Y��L}uT����"�H
()R�A7̠��tw�tJw(J=)�� � �5��м3������`��9w�}�>����}�T2j͡Wf�\X����v2����1v:˥��y��F��\��䢒��#Th�)���a��F���:�������RX֪�$I�y����@���jB������YU�0q&��'%n,�&O�[�qm��YE}�:JUdX��*�|[z��k.�uk�0\�����"�x[���5�0tR#��CW�j�ʭ菊�	��t�'!pMdɭS3'}e�L����a�_~�v���O��ߠI�Y_.��z�i��������f�%���V���pw���:���Ҭ��u,Z�F�Ӹ�|��Y��!���60�L=Z{r(��ߒ�/��67��n=�x�V��4��e�+L��^���7�ݭ���A�o�F$�a�e�|�b�����28����m��>�榬�Qgǿ�Ԉ��Y Z�	�/��H�dE���dG��Չf>�Gc}�\	I�k[�?>�0�c^�R�?�0�%��
Mŝ��F���
;���Z�ɚIW	����]���S[UEw���[�:V{=�A|���f��:H���Ϸeav�XM'����|�3;$E��8j5�t���Q$����l���;-,Oz���(��ߏ+�7yR�_��r��(��=l�ϧ�:c�@ZA9���������b������骛���ֹJ���-�iV�e��k��gk�+�%�oht@��h�S������<�u:�n�q�[�u��߮7o�J���&��W�!�Xٙ��e/��
i�l�Lz��F�W7�y�������
�ឥY���	�_�[�*����5R\�p�f,I�b4�S�C��o��29�b�3�*죪�Ϩ��5n��T��P K]鋫�G/�S�]fb��䡿��gs`��ÏF�5Ė�<F�,�E��mN��� ˽� ��:������v`�]�_��� nR����ǿ ;6���?ΤčVٖ����e{�x\05�1gL�x*��Z�w4��c�m#�96D|hG�:fѲ�k8���mp��#j	D����ԛI�ߡ��EQ�ؘ�i�ո��=��Y���9�moI:�6dI*�ȁ�"O������(���'���Uq��7�/��#s�/�Ф�D�`[!g�肘�*�Ǽ�Y&n�,7�y7���Y��uhh�Ͻ��.������U+��=gF]c%5��|����䣦�ԁ�����x$K�[�6���cZ�Wώ�ל�<-)��|�٪a  +8h����`WD��ݿA��C��[��_�&ؒ�cx@�!���C��5b�/�@kX��Q�*��J}�ﵓ]��f�{���noq�U��;24����U�d��H�E<}���R]�]ޡ3��r]�%�4��^v�����X�Y������9���pr!����rB㫈C`@7�828Z%����y�1���]�2��ܙ��ӧ8��h�����	փOl�O��a��0�������I�g{�p���}	��V1���Cmƶ0�`�u��+�ž���]@MP���;�XO�\~���'�X�n�R����l����' i��^^�#�^�a�ZX"���	f# N��}��*!�X]}|t�"�z�*��f�N��1
]8�����FZ��/� ֨��`@t��A��������b|��HxL	n�S�Vd��e�%%%��t)B���en���/�F��=�4��'�f��A�#|Gw�i��(L|�~r֩}���N�5������槑�9�G�7�F���)>g��O��u[@I�k�7-���x��i�q��x����=�D]4mZE�����C�.�=���4L+�a���9
�6�P���W+�k���BEmDM���X�ؕpx�O��J{S+|LÎ��n���t)e����Yx��s�Rٲ��-���u���G�<T��Gއ�/��[�o�լҍ��1�u�o�2j�d��;�]?��t��k�H+�J'�z���B�0k��u�9��{Ew+3�b��3�m��I^O����@/;�ܶgl�!>�H�磔K��I�A^�(7��jQ�!;�&0���i�a�Z
m�nǅ�Zl��o`�Dg�f������p�z�U�"�O�k��%��Yg&[	b��٪a�����}T���ly'=��2�G�.��z�)�ߑ�1:+`|��tf��B؏m���ڣ#l'��&���l���A�,f"f���#�Uq�[�� \n��4�S�ssM>p��~BG�Py���Y�W~���\D���$����aQ�>�:L��(u.~.�N@������Tzr��<㋕�U{ʕ`ԧ�|?0��t~/��.Ռ:� 	��y�k��Z,��Z��w��D�0N��s)�=iB[.�S���J��1�V�sS�j��׊I��ϛ�!�[6��вz@�����&���7������� n[|���F�����6?��cG<_���Z'���6�(�^ǑD<�j�X�-|3
8����G�^\l"���w����_]���5]�Ȣ�!�c��|�$Jq�>%i��5��%7Eǝ15J��:i��$V= B�~���Hi��� l8��Yny&	w�e�΍'c�!�=�^&?B�"�mw�33�����i��s��g���%�2<�Wj�Z`u~���'�+D��-�q�4?��X��)�I���E-��i|�S%��+�r��`qs�P�vk} �J:�n��k�����[[�/��w�)�����9p�M�n��L�����2��WSl=	.~����&�(���>K[#�SO���]�q�<���L1	^rzg�"�țV|�Ӱ��#��'e�ʑ�?�K��u�a�ͤLҦ�8�7�����J���X�t��d0ʢT?�q�_$Ӊ��Kx�bRw��� ���&�N���G��tMW�<�5��U�;P��)F����b�*>&���il�cV2s���L;0��n�d%Qm�r������@�M��η,�4q��B�_~g�^\�	f��x�V���*�p�$���ʎ��Aq������/a�:�x׈gmEƔP���5�| Շs�̈Z$���zM	?�}y짧e�n���n�� ���HB��׹c^�]�*I�h5�.g[�Bwه��gu.��ivT����d<�0-�/�VuU ��C�?^����=?�'����'�[�����M�ͫ+������̒��{�nN�*A&��'������_�<s�l�}�K�M@A��o ���~�J��e�qB����^��=��y��M��ViB֝k�A���4��_���GS7�e円��<�>�>��{� !~1�H�`�_�(P�а9Υ�ٙ�9��t�J����n����B��è�o�TU��cu��Рgs���7]�QP�Q�訿�-���}g�����|�pSw�[W'�k-.�����I�瞦�.��G +�p�A�. �����}�oޛ �K�R�&���y<�����0kk��[/�D�*	-B@��0���>5�du���$�S~��/�*o��/5g�[�G��BhЭ�h�0�YJ?�tȲ����a�� ��U1qz0���D�$w�����<����.�]2Fy���_ZT�t�t�Au�Bg��oMS�q�������y��7���Zx��z�@��������νd�(�̼�pԢ�I�N�@��R���ɹّ���2�z�1w�2F�1z� �����	(M(���t�h=$�J�N�n�nad~�O����%h�����f7�B�ciQ�y}�adEr0��b��1]�؋�����D|�{[��$���*U6�rs��\#M�BA2C�c�o�\V:v�m�ў&IJJ�� zܔv`Z��j���;�y~��:H�S�ȍ8)=�n�5�q8&4�s��Y�?|w�+K�����ϝ*�V
���:�I�ѡa��F��'��%Z�"��,YY $Ȼ�'r�6�(�G��B���)�f�zv_Jό���w;�������F��%�ЗB�.-2���kNCQ��q
�_	'U���UA77O����8>TyOm�*���S֗��jA�P��-0��Z�F����QNH����\�ék��~��D��6��S��~ܳ�H�����0�p�,@��]$!y�O���R^��%�X3Et�X�l��XԞ��^9͞P*.��o����6o���<iR�4����o}�密2���1�B �-o��|үыjHb��A�T����c��]/�Y!��op�4��rE	k�I���\Ć�2S`���D5����$/��'����/�B�{M>����B����g�W$z�l
BD$8�1�:�Z�=��o���l�u�P��f��!9:�q���?_u���B-�mΛ��L|I�ܠo>��( �����4*���&TZ>�K��4�My�Īc��g�ʻ�xJ$~a������C������aBD�`כs��N���B��L2�y{VIT�,����t������eG�	JV#9
*�a�hG=�*��!�j�qs������-�!ۓ�wH�|wO�
5,Zd�6
&0~����ʅ�S
\��9_�?�&X������<w��uKM�6ۃ�=g��7j��ҝ�M$ 4V�4�F�D���[���Q�6t��'���\W�����;j����ѐ��wc�پP�׾O�8��MB#��J��f�j�j5dy�G��9˝f�س[��=��rݝ��HY�E�rt~��5�J���*1?G4_:*����������p���<��,�ou��Y��*\ �4!"vp�W��&��8#�V��(fm��l=%�~�PK��v����K��D�0{����ie�ת�<���eb����f �H��]��7e���g����GB��h����g�-Iƍ��[T�]�x�@[�R[�W����Sǻ�MoZ�&�7.�����N\�b�êUw�c=�rT��H��o��pKM�$!��ɲ�@��L/�ebv������-z�e� դ�!�J=�{qAq	X}4�Z��O���NDp�?���o�:bj~Ȑw�0��9[A<���fY��dY4�Ӕ#�zb��P�ypV�y�#a�̏��J��x��;����?k��I��R?/���ލ�POc��2T��=�&���9�)j<�1;�tj ��N�?���/�X�t?LR�y��7C_c������z�ʹp��L�ʌ�Ț������~�����C3ϺCe\ˁ`sn%u�xL�n�����Dx�fQ�};p��k��K�j������)1u��E[�����;��)��Zx����^�<�ѐ��E�kv+=S�q���d1�=a�ng�28�0�����	���8��>5���a�&�qL�.��7ޟpӵP(��3ӥ?+T<W�B��6)x9u��H�CK���°�u�6ܽ	��z�����+5�����>*[�ʾ��
���%��g1���y��s��%U�����<��Q�V��(�{~6wx��dόώ2��^[&s����C�Ky,��|p�����7?,Rˬ�g<m�gF��������n)�9h%�� q��_nU�66y���� �U�޻��е��93|��]>�A6O1͎�n�9e�Q��ez<އ��OE��3�kAXXT�o�2��9�~�OǸJ��W�{oy�N�KSML�!؉b=}��S���KE���џ��@�gȚR=n@�x�����]��{�{Κ��A,�>�&s��� ��O�7;�}��\����<��,��ȉ����D�j��9�x㣧��i����h\�����u"a��� �(��V��R�������1�.n�� @c�}?c���H����@ �������(�l>B��bPq��lg�툱+�8�����)K�R=�'9��K߅���wZ�B���T����J�>�xy71"��w11̂�7>�~$^_��j�BG4w��3��*RE�|ӈ�
���>�χH��b���^�Ւh��`��M�PQh���@�]ԗ��G�p5�p	�$y�D����sx75�P�(9!s�:P�|N%j;�@��|��,Dx�Ӏl��u~L�?�p�T�3Y���/V
��q����뾝X�Ϋ��exϸY�� �R'aQ�;;�Bl�&���g���6��,�۞�TSB���G�:wE=��i�����,�`ؐ�T,�#ۯ{�8���d����\>���ج�Up�b��>�ي��ؾ�)�38�w~V�GM,Q�=���S�.��um�Xvi_~�;`y�R����x@>�z---�!L����9��:@&W���r������O�i����t��Yg���E�AC���RNyN�.���Z�lY�][��aZE�!V��2$R2fJ���2�%��yC�
J����w]���sEP(	
Ձ�ɻb�J�a�q��zP���-Ň|��� ��;��Ѻ*�"�^���Fk���f� 
d��	�z9s�F(�\\\�"����PBv1(�=i���<�[['���h��X?!�`�a�<�nXn�?�+��gI�ob�ɲ�	Lg�Y6�����k��s�N7���6sc������+�v^n��!��"�������K�����F���	�����H.,$us�'���$��y-�$9��z/���t�u��e�K��,2�GZb�jn�_5���sRF�?X�ϟ����fR�;�*�L8�_Г>�w�\����ͩRx�pM��)��0h���]�<Y�B�N)0e>�� �sq�Cn&���b��9j�k�9���&,ӓŶu���#�?�Z�?)��P�+K�w�j�v����|�Y�Uk���:	��A4�]���2r(g� ���~�1;˩����)z�p�N̅�U4�=|��#�Ȍ�V��9)K.Ki�o�j��bS�����)��-���و��ʉk��lnŮ�[p.���)�T��ц:@���O��]@c��Y����������V�]*��-��8�)�Tio��K\�0���!�������}E��w��=�j"�W]�������?�<�y�(G�S})���9��6�&>Z\������&��J{=be\s����:Gs�X'{�F�^Nϥ���\�V�~=g<��w��}�����]��	F�Z�(Jם��"�c8)��w�Gq�.��۷fmEOWH\��5��<Dx��K���id�i�`v0ȐH~�����?��^k�fu?;�������5��;z�9��b��\����Ms�w��;N����Q���F���Z7�Nm1.�88m��E��ǭ�p� ��z\?N��csmqX��<���pԬG7�.
?��3�3�!/gý��F�)6<�B,����:�:�%���6��4;o~�q{۵|�����='�]e.�����[/B���F�����+�7�W����D��8z~��P�<"F�{r�E�L�^���?��,�"B[V��M���k{�Q|_v>�4�=Y
ן��K_2���G���⠹�����}�$�<�9NgrҜ>�|*[�8ⱗ���\����h��Y󉵰�BK{,�z
���\�����{X7�z�A��9G�-wU�)zF�֪����[���VG��n}�efu�Ё�;(��B��!r׹-���հ�\��s�+:!�,�*V��Z�N%����qxo
�hJ4�����z���L.���8]juGM��ŮL��Le�y;� O'J����~\�-�y҄�*kZ��XsXY�g���=��_dJ��i�E
�������<��6�r����r��T7xQPNFf�Ƕx��k�y|�~\>�{�%�}��9r���}t���V�413�;�Vvo/;��Ȉ|�	vV���Dma�	?�,�-pk��3)**�\�Wr�I�#U܋�{�Y0�GQ�K[[[?�>I�������j�Uk�m|�`��#ח�f ��q��]�ⶦ	��Z����t��_�IJ���#z����J�۶Y���� ���%w	0X[q��ȄSF��ԳW�"��x�'�
v���������{�w�4�x�t���Z+猴ܳF�}cw{r<�V�*3��`�h8����W��ӵh���sW�k�-��M=���Zv�+$�NR����j�rA�	Loc��
�Ə����(�;����D}���3k�Y�
kMp1�NY=llB^Sy�Ū4�en�E)���A��Ҩ�}�	q�kY���E��N]Lk�X�l$s�.<8::��(����=���K�C�������q��tT9M�"�*��1aĈ���G1/.|�cɩ&��kcm�[�X5�F���7p��+��\��t����7:oȟS�?T]n���'
(y����5�d4����ܖ��C�y���g�%��Gh� 6�2,k��۳����)��nذSF��K�x��,��H��\�� �.�l{�	��p���H�R�~n�����rlIRNG1h�7�sb�+��uH{���I��v� �de�`T���j�6n�����Ȥ��7_�܆4oA;Nw9���Wz܄��g�ٚK�Ӽ���y�Bu���e�$G�^4.�"��."b�%B��:������S�ݯIVs̽�iim�Ĝ��bBk�"[��O�1��o1�I�{�����aHwq��s|��-sG@�3�e����cL�����Q��05��u���N��.#P���3:{�����L<*����2zhХ߼N��!�F���\����x]����ɇ�|�A��Lm����cqB�V��bd�є�<$����$m�I���d?'����&���"j���`��1����OQ�K�`��\���%��M����s4���Ǥ���4Vc�ǵ--���r�+�Q�z��d���wA`�Ne@(�7ȑѡ���(۟%u������KZ'����Z~f��R��较B�x�s}�c�s�k�"wj7�J_Ǧ���.��/�kI��STId&|���9��u�J���f��\B�T���v�J�DAþ�yƤ��j� N&�ŝ�^j��NO��p�(w�{���tَ3^RCx!�������U��t� ���q�'�X �2p$���~��ӆhU�R��Ɛ*�O�efZ�t�W����i�4꨼=i��b��@k8�E"?���=<�*o$�N4��n{s��Q�mM���K����v�ræh����d3U��.�J�Y��A �aB�/�;�9t*�c��էMLW_���Z�@��n�95!*r��D]mm�|L:8�h��V�o�������-��~h���$�V�}���͌ڄ������ח!A%Y�1qH��"��rЫ��gl��S��Rp'���8FhI_ɍ����#���H����Y�׋���8�L0&��q��G�B���u�L�D���u(�������5~���7V*N{<���*I����8)J��4�r?ܶ�bL�IEY�W��woV�����]\Ȋf:E{8B���,8&D���݃�7�,��D����o�~����)u[.�)�c�M��4�K��"zB����:H�4YЋ4ϲ`N�����t����ͯݖ~*�z�<b��5�J��ɖ6��-��/RA��,��g��tw��d���o���S�L{e��������]��ZIp�<�&u�r[���Z��y�ڿϘ�
&�~��Q� ���.�۝2B�{�\��� ֖G��%u~��@�lrÞ���XI���×&qbP-��A��������V�(��[ac��p�+�"�ֱ$X�.�+>���)60�r�c����j�V�l{�Ԋ�$ ��<>�q�s#��:� �ͬ=�!����m�8���c�߬��_���?�t�#��j���~a����^��гB��;�i��v��?z�x#�ECM³syL���m%�C^��u��B�?���O>���Ů	W��0��n�E�wH��_f�t��
���.��>C�6���M^9dW�b�L�Ѭl��F���<N�܃�(�El�'bca?��a#	�"^5M�8ڥ�����8_�nv��E���!���7���l3����kK]�q���y Jje!��f�/���=����u�Y��"���#�F(ϲN��g�``�FX�"�A���|��孖��J�v���0�I��B��i���'}x�gX��E���h4ѡ�j�E���4o�O�rz��{�������@���r�3Q�)5Q m�ʊE�W�{3�V��[0Gq��0ԕ�a�R��̓
N����q';R�U�~g쫃C6f�GHG;��(�����Q�~W�.)�p����?_h�O~���E���`�3��ˎ���Q~1x��=~����$HLg#��zܞ��]�F�q������h����tꤨ"���^!2�7M�%1$�Y�Fʔ2š�����z��s��uB�}���6��qf�o�����:IDt��D�x��l��2_"���FV��*�����7�o��z�d�d_���j.�d���I$���"���?��J&�]����ڲ���uXGJ��j}��:&�ydV��6�QuM���Gx��BC�=l��(���-��hS��2���9�yD�̆�6I�͚�4���| ��P�ըOW�D�5��ߕ��OT	���Q�]�GW�悒�N�0�^hŽ���9����^�'!�������B�~oV[n���?g��*><��q~gE��ҥ�1{�WW�T�<�@+��ot�
�|��I2G[��Z���d�Li	G���c�:
'
3';���Z�$�>x�V�;�����| ����\h��lڞ�6D�9����R�����=ȎS77��e�jq2�Of��p��ޯ���;�d���o4}���K���G"�M�3.�{�a����=z�����F��}����8I������j�h�Ar䍻�����KS�Ompk���W��Ï��D6[�%ade���Q_���lZu1��E���]�l�����w��
��a1��؜C{k;�v���J}��Y��_ǡX�ѯw�$�����d�ū��B��g{��J|ۀ0���o�}QϜi3���Jo��a��!N��r�JD�DKR�|����V���Bq�D�Yֳ�jɚ'>����	iY��K�R0X����d��~|R�+��ڿO�%|��s���}ٚ=��y� �?��G�c�i������X�(M�p�e�f.{ؗ��(�ٰt��><_���]1,!0(����� �X��ٓA����?�Ur�=O������Wz5�nz�z.�@��v�5�]!�a	˗4��N�2��)JN��RO]TdO~�>\�A|�so�����4��Mq��,^��]8�>΢�f�����ǂ�$��s�E|�zm'�0�S�]4��g��7��@������l�K�ċt�'�v��ݶrd#��j.J��a�bv7���+��sr8��	u�����ڸ���1���y~@U����\6'ɏ�� ����Cw�s���0��5S�K�(yv�o�ML�}j)����e��+UAn�맫�ǜM�+[F��!;k������6*؟�`�p��B�L��*W��+�&��p�ϯ_�C�*����Tq��ClMt��-e�kϤS��1\T[fwgtu�c�GH�"�J�(:�C7���T��W${$�y���h���A(k�h�rB﮶f�A���矍Q�¨O%�a�1sa���`���c����?�um>��9\��;E��J��*�Ԅ�2� a٦��)R�'
k$v����e/��u��62r�"��P�:�Vs�	�FG$2QQ�Y�i�yr�BU$E:!��Q|f���:]|����s��f�����q���}�u|����,C������}zU�s	�\��9��m/J|*�����j��(6|���e�_�����Q��U�ϸ1O������_��Z�t�M����7��X"+�CR����s7�c,|�t�*�"�^���ǽ��X�K��l{�|8W���i�`��?6�rP6�u�c�6C-�?���7�.��υ!C��vm��	�B9sp�Z�b�q�'��� �����!�+�ytH;|l��*���һ�4)�N�w�ӱR'	����[���(ɛ�����z�K�O��?�@�`�t����'����>U�Sy]8{�ˍ�X@Y�]��ׇTmΰڊ�/�ܝE�y<s�Fv��c�=���)��- ^��9�b�e�� Y;��3�u�?u����|�(1s��<]t��Yg��_�i�O�]KV�,��"��7*d�5�?�o�Z�"C�{Mf�+�US��٧dh:��(ج����XA>����,�7���م�?TeN�I�G;_*!@\QKi,؇-7�l���w��ͦ��q�[H��u�P)��Y� �d�d�� �0�L�=�d�Ȟ��m�8�����r���~b���!!2���=������_�+!�g���oy�92~})����M��<�^F/�b.37������	������9�a����#Ł� m��Ϊ�(�E�8D\�S�U.��*����mۘ��т��N�$u�����ع3�y�P6@���)��om��ϫS�d���Hѕ�8�W��T����u��q�iw�U�QD�u-g������!�໷'&�����$t�g�~�r�l`S��w�f$�p
J3�F�g�녀�H�c�G������v^{���-n����rm`�������t��)s�쬎��xAL&��a�N���0>��̯������p���nVgK�t��%#D���Ƿ^_v����h�����/�J-�s���#�|r��X�{w����.��1��͟�h�W��z���e�d��M૸��]�uc�
�ɔ��Vp��u���֒���ЧJ�eɳ�h�������'���u;�0����Q�V���ΰ��	J�a[w������u��<ʱ�Sq�ʩ��(4"+����wg�DRl����U�`�;e���k�{���x�l�{�I���I'듨q;3_��7����鱒��4�(���j������!{=������%s`��KTug��-�{Rњ(�����p�=�����K�pX���j�qWA������&��Џ��Ct֫�~������h�<�s��9� �H�H.cnV��>.!� � {	7ec,Ó���al@�3'��R܉�;��������E,�b!"��X�ɛ���\-�o�j��Z������=<J���I] y����!YcG����9Ӳ_�ON�a [>V�X�L���+!��=�	�(U�:�p0�;CW�Ҫ��mz����V�n�(�7&����v���{Q����u�D�1�Cs���w��(O�C�c�^A�չ����?��;+7w�\�7oBE���\)�D��2%�s��n�5�A1�l��:
YZxA���c�Ղ<��7���ڊ�w��C�T�5����v^'�d�+l�]%O�sS��ս�P�ި90J����طB�N,�h�vɳ��K��L0�<�~u�>��y_@ό�5��$�����%���+4]�Ⱦ�݃R!��F���Ӿ�\�wD������6�����]�/�����17d�E� u������s����Ƀ���Ҽ�읍rJU�H"����1r+�ą(�8d���m������c$��͖+����D�¾��R�T�2����[�u݆+�LN�H�L��Jr�W�y�+���>&�gVZ}%?�>�z�\Dn`�N�2����!��A#��3���G����\�q�/��v�J�J�p������zȶ���u'�i�������Q��a�������j�z�u��}'�J]��l����[
YZr{m�+�]�h4r3U6ڱw2y�vny���	�Ő��X7֌p�<�����o�!{�r�tn��9X�`5���Qkv&)Y�����XA��: y?�A�o�,�,�3y7��1tE(�U\OM�E�[A�^
n,�����M�K�(>�P�Fz���Z�鋮y͏��5Lǘ�Z�8���T)7Y����O}%����F�60�_�3���V9��skS����g�m�D37f�-qmB��"ĆZ��_���.��"z����%랥Yi�.��^Ail�a����F}��իv���\;1v�e��L��o�!����Q��v��y��d筕�7�z?~y��&<|�{������Mw0��	$����M���Ȯj`_믁��FA�k�����3t�OA���e�(�w�;]y�Ӕ��c��{`692}���D]� J��,	 �DX˹3�f���9��N{f`�䌾>��-�������F�Ǒۻͧ)�{-±Q �����Z;+��rW����o�g�R��Nv���s� ��YK��A��w�*׫�����D?6��S�H��{��{�%d{+;��z9��m�t��U�jd��������-��K2'�����ٚ�p-]�nİ�����.C��㸯�6<�_=3�?O��Z���ע��ڕ*Œ�
=ht��r�-�m�w�p}�p��z-�p�CWeJ�j�B�����d`����ܓ��:qC]ݟ3[�����X�e4�o�oG^_ӓ�� ��s1-xݰӐ:pxprJ�� R�0�F��*%�q{�{�S�����uh}g�Zn��{g�O>6�hiߓ/��~�0\!�96c}i�������*�	�LW���t�?B�z��;q�Ĉ��~݀��\|4%�5���Y:�vԧ��s�Β�E���^��U�[ݐs,���>���v��@aY03@e��4U/�y��j��jb ��r&_�o�~v���|���*`�᪖�}��BV5�ǤK@�+��k�����58' � �9����d��pF8)�_�_'_�Zε��-�A����s�Ng��^b�O��Ԙ��^o__���lM�4\ː���M�D{��5��z��L�Z��^�����n]�O�{�}��`o�L$����5�`�W����E�H�G�?��z	e����|�(�h��	����(>cuG�HoQd?�A�����n�+���\C������������v��n���Y`�۟f���W�ep�'�RÒ�
j��>j�{b���f 
�U���N�Sb���Q<�T���@�k���F�QƧo�/�;��z�Q[P��j�&�>6ӽ	�A+��e]@O.N�h��` 
y����������p�� �ba6����%�ݔ��4��/E�ޚ�
�z��"���5���WjL2�˛ϊ��d5��\Dx��˂��a��1G�B{������T�H��j<��0�8D���4C��@�Ã�/���9�쥯��1����z�����q�%#�m���̜g\��:İʦVQӛ���w�*�%�	�Ś��ry yS�J��xD[J�^���Z����Kv��n���"�[=*�;��Sc�W����k9���~K��^�0k�O��ռ���1'��1�ҟ��Ő�J׬�l��k�ix�=:8�ŏ�_y|��&E�L,����(i]Ŝ�kߖ�䥩�ܶ�6s������;�� ���x�0��/������y��B�l����:�ɆQ=�Ō�f0w���,wm�"�r�)r�ss�KU%����!U�?�����_���zQR�L0�v�s{w�uڻ�%����������]D�jY��5m���Q�/�^�D�����(��>��S��ˠC��:V��]��e0m�,Y24R�#�㔉b��F�����h�G�yO
RD)����1�^��ॕ���k��.ׯm}���H����_�/"bQxm�JMIᗒ�nk�c���446q'L��1Ȓ��FΫ4�`��j1����+�S���Oa�L�M���P�Q���/���0�������R-U.!j���/E2����{�x�5%�`f3S܄��u��L���͛�<t��ggg�|���4V���]�t5T��!�k�A�νϝMv��u_)v��^���~>goP!܁JYu�(�)����[@=7�~�;f�s>��bv$��}��Ȕz�?�^�G|���#lT����X������1!b�U)D��ƛ݆�hE�0$�>�X�4Q\y�x�\���Y������ޜ0sC^(<(��˲~�n�FS��S��G+O�4;�{E�E���Y׃���"R�Y�ec����`��_�K�fu��Z�H�)R=�s�M������#����r��U�]3\sv�秳��z��إ
���-T�-���~��� 5L��[�o��/�����<�I�OGd���(�].xܺy?F��;��m�02�G��-�oaoA�Ӂ���w�ߍ�+#�n�����-"���]M��&|��!ZvhR�
[.^r'���N��Қ�����Qi� �^�������s��Wt}h9�Ӷ6�k�� <�#��3ٸh��������%�}5d LR�q���������r��o}*��W,\��:q�?�vK�$j�3v�9����"Q��_#�|a!��t��9��
�U{��_TT���,��~b�7���ˆ.;3����:h$�B�����tb>ӭv��vfS3��C2�P!�!���XqK��r:��7-Q[�/o9*�"w��ܝ3b'5R�����K�cm�5���9�_��:˄ֈӃu�3��u��~d&�rl|�`�b����Z��mKrwM�d��F,����mί�:�Z��-*�c������=O��ҟl��n5G&���k�O�i0ƕگo�R�����j]�fn��+�D�`��D��O�7��No�j�>�Mi���c��~���P�,{$�$G�Ǌ��lG�
��������Q�&78{�P�q��͝��{_���~���ǽ_���9^����K��k�r�R� 4F@�
�q�c6���e��j���`@�A��/�d Y�㈆�4x
�'_f�����+��ѷ��R���ܑԢr�Z-.���6ǻZ�w^j�+|�bjsg�I�� +"��٠1qgh~Y_$��w��=�lj>:#x�i�3����p�����
a=r����awF�!P�٢��Bi+��x�bd�z#`B�\t�X��U&?:m��djju�"�t�w��Uϭ� B������S�OvF���rNk+/oA,��o�7{�AU��v=F�)٘8>)��Wy�'"���W��eQ���6�堜&0��("����k�'�^=����m��^N�`�5��t.�ez�0}� �:�1�:��vM��q�`l?�z�3&���b
z27;�U�~�"t������wL7�	?c5��h�Ey�5���]�5�ps�q�[C�7�z-88�{@`��N��()��F,qᛰ_p�&�f��t����F?p�)۬�v^��%N�
.*���@=%���<��b[�C��w���(��[Q����ۃ{��8����5�nL}����ks��ppt[�U&�߇"BF�O:vUPg�	����m}
�=xx
��M߹���Y�0�{�]w�����'�@�xi%��^���3�>G��m[�\��6���������xT8cUd5"0)���OS�P��`OvΎ�����ي�56O��|x���9�Q��+bW��.�c�Z}����Ib���N۞��牄�y�U�RW�D���Ү�-�L��ɺ�67&	�
BwM��f�P�K#;�K#^T�.ff橄�׎yE���m붌���L�L�sH��;���Ҫ�G|�K��\���kB�M��j��/� �c%��͡���|�Z|�c�f�G�e)�<��p�������� ���[�%�r ��&��K|�tPI:�j9��}w�7���kH�{������ĕe���8AO��%}��x:�DRR�g��v��K�e��%4v-������(4>z\�#���r�bp���q���?�?2��cʭ;w�K�t���p>:F���ɪ)��4aq��G�D�/"JEg�F�5�`1O��u����2ɼh�\v���9_��
jw�,d\q�U�n��;� ˙)��CL��ΜivKл~����(�2x{,�<c�r�de�c����|��K?�M�f�S�l!����I�����х���_�U��N��~\)N0*e/#�}G���}���]�"Y�u��5�rR\�	l�u�ǡN�j?�5ߛę �`cs��U���xK���3�h���)/B&H��昂&A�NU�	��z�6��)��Y���X���JF��N�_*��Av%??���_1A�ߺkP�X�Y�]�*ZhR=����;�|S��EsƢ�8[���]�hp3�̯��f8S�Z'CW~��X`����fDF�����y��:?�#y�^�L�F�L�ɒ�~B���?�<����m�3Xkc�]6x�}v��' �:L�q�,�M7��^�*±�����)�mb�A��W
ȹ��0�(����Oޗ#��s�J������#Z�`z���A;�<6~�)F�*��ڜ�����$� �v���L/Ek�!e�Ҩ.{��ٷq_�B����	qa)|6�`ft�:iO�}�'%~>���� E����ű3�+���<����WY@��O�>��6.�Oz�7�H_��}��^��{�w[$����ڟ^�Vq�u��_�I�R�DF���kE��CQh|�����QL܃���(c>�B	s���+������ ^����܇Z��~�~4���S{`�E�(�#*t�Q��ʢ���^&�y���d#��El<
�i��xG�/�Z�0&b�_{�����U�1���h;�#&m{J-�Aޟ�,�M£�C��J.Z�1Ny
�8s��$5՞�@ϲ�]˅T������Ś�����(�V�ᜮOw������s`����|�n|~��7�`�8����cR���U����^j0_Z�TRZ��un����H�
���S��҆�k�)xa}H?OZ����f*��67 �ޙ.�B{y��x��r���:Ϗ>p`�!��:o�L��:����*QK�w�h�����[�_-q��U�!�HR�W� ��C�0޽�3���?�xN�4��.�����35�� 32�Ѝ��O�8�)�$NGV�\@�5����U������5�^�k����,��ٷ��~ʘ�5J[/��27&0��ǥ2��ON�+X��g=92B"¾s褂(�>^`�r��*Z���ǚ�|������$�ӨL�K%𶼾B���"�U�.�3�b4��tKw�Z�N�򭩈?������<�v�4���`���qm�Qz�\��z�����w�6kc����z;y���L�-���.��'KL�Ψ�8f��Y��Z�k��*6��������.����;��AmRW�3/58��O���q��$���V��&1q
$iM�W2�R0��V��1
���,>@��Z�s����g�/��E�·�*���=J(g?���#=b���)VJ����ˈ�z�nP��;��zqO�����U�������z����_(��1�٭�_�:O������?��t�3(�PB��.�?�@T�HD�&2c��R䂞R�*|~&�)��*h�\����߽�<�<"6T�����[}6M�E�`g����:`ܱg��9�ò�,�m7��ŔlP����u~7]$��L�<,����3!�BSZ���0r6�5�)�L7H�!:T��������gTA�P���CËY:�_
�Ҏ������x]�����,��)�/���WN~+~�+�$7�&�wvH$d)�̍�^�^��U�b]��&�p+����b��j]�v_S�,��=������"�K+����H�{<�l�ȳ��2�GS|ɫG�E��ڦ�k�nP���YlL����c%��޻TO�2����U �������J&�x�q���4;;c'���m�U?0�	�?A/m,���
'����
&æF�^��K���,���I��˅9|�#ٰm՗xȉ�=�J\�4�V�h���)�u�|�o��q�0��W��K���ޕ?Ыҷ�v�5�թj�u� c�b�6��^��_6��>�떨he�/Q��u��20:��.؟�[���o��qx�T���uP�#vǯt�Urs�B��X�n������<|��g��V���z���jp����/�� ��"� �͉_�Z�����H\���=U)#P����~Y��>��ű��n.m��i������c~aP�>T~�����"&D$C	hM�gS-	��%WG;��t�z����<K��*����y��������~4ӿ�W0���\B9��u�Wv�JDH���.n%�f)Bq�pw5�+��[�!��I�^�/�v$�o�ؒ��	�&ؤ�lT�C�8-��^�{`f�v��p�\��i4�d��z���\�d�����rt0�:/s�����!nY�G~���OJ��@ Y���{���L,>�b4+�������X�%b���>1�rD����%Te�ٽ������{
445模��/�C��L��R<��,*��)�%�u�%p�%�b�����:����A�I knOxnv+W�ݠ�<��;		r���v�ZdLV'i}n;�e���V����[$�F��Jˎ�l�q��e�LH`E����b���W,�x'L��[Ak�xy:����Z��n�⋾��Wz��f*�!�f)��t�c�����ܫ*9ε�]gˤf25ă�c��h/mK�{<�{��'��9�Z��:�9�:^{�솿0�$'MCIi���G��|&�8s���b>����l�޿�4�*#XJ��0���\uF#��=�[.�ӼW����ٜ�_y���c!0	��:��&��C�f����4�_:�����R�Q�!/0|&~��j�^ �K\z(��Ԓ���E)9E�?~3���*QK�P�E�.�3�/�2��`8��-�#9E�Kz~�g�� iIڮ�f��-��Wb
�uS�vj�
�XkO�X'ݻ����?�#��	 ���2=NN>c�Ab���~�_i,qbRe�e"J;V��d�J���e�.�o���ުI��7S�c�h443)��r++�u��&�p�ґf�5fJ-
w��KCo�AA2���0���t,y�z��t~Mn�\��ӽ���g�E��LGW@��e��۴�	CM�Z4�����&��~i��.��4�3֦�����86�X,�=9/zC	�^��<���2U�O���i�Ğ �����IX�^��]������l���M�E�~�h����G�ZP�T�׬����L(X*H��mQr5w��J�P���\H4�7����1N����L4�\���k�F�0����:�s�W��,��k�?�f��J7�П�Td���D�0�'��^A��2����w?���n�t1x%�VѶ`V���~�ʕ�{،�TTUZ�ku��g����E_�2�Ӹ{�C*�+I}����J#��ϑ����ɇD�*a�wp�>��q;=+�6��PSU� �{��L��M�a��'6�[y�T)�.�}�%N����)��(���A�4���[zf|���໘�A��7M�$��*��:8���y�*�%���uXu�WOȻ81�%'C#�Z�m��u�����~�]�p��
.J�S,⳵�U҅<Cb2Q��������bn٣��Ɵ��:6�9i�3e�S'�CDYbM��S9S�����1���I��وG�&[�V+�B�?�����A��pgB�v�>�Gƴ�Q�BnΚ0p����E�2��I������X �1m������adG��	��i�!��~�f\Ԭ��w����g}	?~z��]�8r^q5"��S������H���+�}�)�K�g�ӯG��M�W�Y�
�L�~p�}�j�;�U���(�7�\�C`�->˾��w���ƻ�`��o�E�i[t��D���P��Q[�7ӭ�$R�T-�g"PDm��$0�Ǐ}�R|z��W,�'ф��%=�$�rZ���6�B�d�G�ezQ��n�҇�>ɚ1נ���A����x����&�3�1�ͮ�y�%���n��u�Fw͔�rt�3[GRɄ��Y?�@����ٓ0�}\�d&��j�S6:0y��/�]��6����l�;�E<DוM��s,�O��(3���v��<O�����<`��<��mv�\���f�D���,�2�]>������<'��>�gee�x?���8�D[�
�9	;ji �c�<t�B����lUJƚ�R�/����jg���͈MT�!<;g���/@�A�Ģ���<CKɕ�gz8�T�f��IP�}Mbؿa�s���|I%4��Ϧw��Կ-/ȳpGݷ�������s��x�3Kk>�LZ�Ҽ�x�r�@��^���t]J��{v���P������L�P���xX}L�VQ�c'���`�}������3�a��O�����o��'�ՑRJ~í�@L��`�!�(5�B����d(װ��%�H�Zs�ʩS�i�(zL�̲F8�6�$��^�3������LNP{�6)�\�X��P�wF����ȁ���|��d�`��H��2��7��@H����|��8nHПB�|�k���A��� �nl����o�X+�q�*��-lvy)�GJ-�
�l,�r�6�[���S���ZS�z��^!7ЪlO_�ӈ)t��A��/ʞ����_��|$�;j_�F���Րj!��k،CH�H�c�+�r���i�T��P�嫻�c}���
�>iY���Q.t�7�u|��b���#-cp�kTϠn�,������Ծ���I
@�<h����}��go�D�a���kk�d��w6����q�����6�U�+o�FWG�a�]��ۛ��b��0��[2���>	�[�T� Ŀ��?�D�k�YzMV����v�9M�����Bt�𲊊�o�y.l��9g��V��Bg����n�K�%����ӣKŽ"�#>od�����X&o��[�Ք�T�&4��X�8#����/�F\�Hiw��_Hv�>]���������dm��;:B��.����A(eE�_�Z�2���P��xQ���v9W�]Ffk�
�1ͅ3T���(R�O�]#}��n���)�k�-�w��YC\"AK����<_��m��T���xBʥ�ndH���O~d��8qt�Q7����n���[��w�u���X���e�l��zJC�W��V�de��[�=n&$�����msF�O�[-�8]'�碔:�j杍b�g/f��"�4�t�kBc&|0�Z�#NS\���3ӶN�!*�/�9%�ۅ��յ������U��u����Q�e��	����,+r�h%�Z|�L
����e��Z��_ؠ�JT�Ko}wI��7W���		�W��X�Qq��~��Bnd"���s+5�~�0AK�SO���e�!�Bc�'�����Q�#�F"�n�lo�U:Ϙ������H���?�y��q����t!lS�9
q�\N2�?�_YW��$������Z8�����[����^�A�!��~(�f�ؤ$�Ms�2�b�p5�-M�O���-h�Sud��9�-�HX�����+�f�ip���;����;���'Hz2l��ى�K�nݜ�!�3:fO-Fc W�DbZ߷��!�W�m�.{
�ʮMQ.gr����߸������G�;>�(�H��KMO�/����:w�Zg�W�����d��,`����;�ԏ-޽�?p���`�Ǽ�wGGd�c=�?G�G[���������\s��>N��sM�
�U��7S2Q�~hL����w-Ż|�'�^(�n��͢>���VnU�r�H�_0����Z���s�z��Y���HF��'��f�*!Pj��戹Q���B�<������:=��A���Mۘ��������1��Q�p�(W�d�?0)�N}Y7��3ڻh_�,�]1�w/�S�O�1�y+:񼴊�9�ش��.@�m��\*e]����m���.i��@T�}o�DUF莖Y6���vp�H�����B�f�kQ6p4K��ZD,ېm���&,g�<��}�FG���I�O�����[���;����<#t�c\����S�t��hm�:ky��^0W���H�$�ΣΎ�����@�*�������I9J��8,�V���Y(#�_��#�P��~�Qw�Wֽ�-�:�cYgh��h��Hpl���\L^y��B����n��>Ș��$��'��7�8�j't�A���zA�x^$����g6�@����i�e�I�^���q��]��ǫ:c����UI+jQ���m�t���B8�����R������z&y�Z�0�Cjd�V{g�?=��.�q�TkSX���~I�":��]�����4���lUn�v�����~��B�g�̕��5�57�Z�fF7���VTk�3�,tqK��ܸc�}��xS��>��n�}>��H{3�����J���k��Oh��]}��D�d�ݎ�<=D^����D��,�I����<9�<وQ�>U�j�\6n�I��[4����`j�t�O7�ձr�|��j������P�M���ۻ��7���I,��ׯwI��|����2�܎ưX�Kم�o55/��&�� P_�~tTқ�jl�^f_�>�>���ע����S��4~�p�uM�{�+MKP��z��0�>6����^ŷ��{O�&���ϮlQ[�ڹ��ͺ��h���{���%X����^Z�ܨ��SEc�Y����q�Vj���ՌC��/,1e�dD�˙[+U+ˌ�A�����3X���_�ZҤX7��CZo�nD>ŭNp4=��/��UE�� +o��5vr�ן��3�O|irE�nmgNj�.n�z��@��x��S�C������X��)VcΣ��k�mn�jЀi�R�]�T��+&|��h�d��������\u�B<���;�vǬ�LS�K����OhR��~%�u�����'��)���L�����OLd�Ĝ|�_\WB%(��О���.�殛'On�1�>d/~U���:�}��y���	��z���(+֔M7Kǀ���/=W{v)|f���l�&��!���g�Q�q��ɵ��w�5��h���2�0�qb�h�V;��[v���^�w�v�KS��3���	���60��=�$�O���I�w��b<�}�,k��S�L� yUv����#��� ��a/�wV�M��2�`cG:X+�_�������PF����v-��p��Ȼ�N�$N`�n��Q8�;�A������=��\������}�MCC���F��_L▨��β���E� ���!����㎎�Bk$�5��`_�kaaa����@J��ɫ�������`aU?�Z��/���IR�l�k������P��p��{�n���[Ωa������u?�\��G�Jbe���M�z(��*�˖���5��LqeB<�,��/+��٧����	�������L���8$������o��Oq,I�vFu�LB��<�ݲ�@�_e�I��a�U͑���wզ�{��S#��;�캎���>k��o�F������w}�(�>���11μ�8{���
{�e]F��7�ag��X�"ʋ��s?
����_cyn}/����N ��g�Iq�����/����5�^Bl��ޛ׭�b>�ǟ�p�p���U���dMLpQ��JA�=���C�2���U��9�>�$�ײ�ob @g�R6�n�w��,���Խu��v�:�����=#(����7��|e���
�o=���:��I���1�G�#]4cS�y���̀:����+��ѶV��*�rn��i�%�^�[ �AEW��	V��:&^]N�1���l��Xκ�FO��>�V�~�ա77K�Q�,��7���րs���G�����*����1��v��U}s�H����	u��S������RiG��j���$X��LÙ�wD9�s$�?�T�xSj�޺�	K��~�7vav�����~b#��nŌ�u��������K�!���6�׺V#9�o��e��0c�>���']�u���\{l���������B}Y�k�AS��B��F3�ޖ�\)��Ҏ݋[��i��Y�5��=-�G���'Gʯ�9�s�eB�c�FK�K?x��I[N9Z�o7T�d[y���͵*��]9h<�K!���	�?�fF~E�Tp��s�ظ��X���;U\��Sv�7�7��ه���;z(p�KSn�����<�/W�m!w�y?��J�ȼ��v�����<��0�=��������dGњBCㅫ�%=&���:<}R��$N����l0RQv��眿ˏ�^i]��R��t��^�4�]��3	�K��u��)��ąg��y����Q���X	ON�'�w�"�g�:��FWVƐ[����Xb�yQ��ҩ���j�KV��D�ڌ�΅ɭɆڙ�W��6�pZK.��ry�p[�[��*�eLT�n��np��*������µ^���?N��岒�!���%[
�����\�{yC�?��R����L���]��O�U%�Y����g6�.")�aU���m�^��K��F$�����p���������Mc"<O�ɸ��:{�9�*{��w�b�x��<�)╩�����!���(Og�<���aE��]�0JS����%oF�`��o8(Z|u��#ా��6�R�8�LMM��Y���[�mlX����['UoE�5\��=2�e3e���:1v��c�3:�����ks1IC̠�*�8�ޘP2�g�kФ���M�Ԑ��v�t�tRu8��Nlm�n������F����΢��N4#���B͵��~�!:�����f:h�2Qw��|�'������i9;�h[CI�����q��ӈl��}����M�z���H��*��u����H��brn���;�~�����+�̋(���<��4��Dy�qǎd�
��-�u�z;���'_����i%@I��p����T.E�Y_����#/|�G��+ꎫ�.zډ�N��-�-��'�#N�ǆ����}IWt᣸���*������[3ʃfd���«��iae��
t 9�|�	<���ã[��,<���.�.�5����7;�N�]"����<�N�?��V%:^�U��1a܇>�k�� cBr��3jnH����E(��]<�[�°.�J�o�Nxa�r�V�ت򆠡��߰��u��
x��[=�D�'��GGzt� ��>{���<���O8�-Ğٷ��Ϊ�yK�h�Cj��X��7;/n���(��x;L���  ).�kŬ��%[V7��͢q�@�Ѯ�R.�A���kllM��$>N֗�a�G�'��'�����������Rc�Q��)�; \[�l������zK�4�%>t�l]}U���l����5��b�=���H�t�E qg�Ýu��hc��6>ԏ>JD��o�X����8ʨ4�����[�*�D��\����\�B|ڿ+���)Gue���_��Ǘ��9���(g��d��#QW0E�@�{p���m����.e_�?�Ԯ�<̾׎	>*�c��aqy}��$vi���1
��0���V�ޝ�C��ЙO��s��]���LqIm�dۆ�UD�Tu�po�_��dF݄CY���%��{����������ki����Ķܛ�8���m��{V�3b�u�r�N�������zM��dz��$�͠��%JZ򺤅S�� \�m46lK�]���A���&�%��_\���e#�D�n���F���m�~��P�M�)�b1��������&J_���Dr�->oo1�<#.b�q� ���f�E��b�0e�8�\����;�Q*��%O�v�����aS�"o0D� j$s�/�}}B�����Y�	���_�ћ�Ï������}�D�PȐ�i�m�T}����&%4O�!B@�/�{�%�3�D�����
!��� ��0�xf�����	���J8�<�|����NA�+�ؚ��g����Ͻ�����:6�׀�mu�m�j�#�T���;_9�x�����P�-�jh�!����뒻�X�A����I#CY���]�%�B��1UJ4\Z�c���Ո8��"�$��sgy�_h�4��U�&��ϊ��|�P+�����͇\�F<�ے�?��EN�sQJu�t"d��d`�qsrОk������.}�.&�;�&�(*v;_����n�Ϡ��%!7���*3���F$�	ߏ]���29��?��B7��՟}۵�W>���������:�)��eYdy�'�G��Z�Q·������w���ƴZ])
�oݵ�Q�z�6t��oߘbۑ������O�ֿ$��l�-8�{_eo���vx|�(kM	��'�]�\0�ǍjL$%���]��T�cQ6NF����\+�w�-g�x�_r��`�fG��l��߆n�'dU&�a��ٽZciI�J���Jۂ�Ș>�]�C���t)^��sjs/��"M$�5�(Ux/ɱq\S+XELMP�n�|9m.�\����-�f�+ rw)7�z�;[Dd$tu�T�6�/��Wڇ�(��i0(X��|����/b�a�g�Ӥ�^����U�G���L:z��ç^�>���3k0����
�� ���%��F����!
M�?FЏ���+�/ɫE�ql�<��4�o� :�2n�W��H$\xX>T{���˼ǿ{`�>40����\�fD����HL��<��=�sz(���MK!�s���vaycK�f�.�据�S��
�{����hm��Hܺt��]Ϥɿa��@�(���Ӆf�Z���ǭ2n
j~�;#q�$���D�}<�{g]�"j�r?K�`�x�~8���"�\����
��bL������w�������x�L^l`����nc7��|/����>�\�܌�K/t�W���W2�x����ݬ2%P����1��&�P��˷-�cy���ê��&a��"�lO�Ѯr�m�Ye�-�HTR;̝����0�k��eC�|��҈�q��<��P��p�������a)����=�����\��5gW;��I�x��oPo{�|�U:?��I��=0��}�ECp�b��u�bɀ3�&Y���;��z�������xN���O����OpD<���P�|�9�I3+��4b���j�[��%�8#R��%�  C�,Qn*~�AvMM�RRU���^^2�u�9񎆄�	q��/j�#��EQ�o��:��SA~[��1�Tt\Z8�i�J�Ã�+jjs��Y{��c�W0�r�Z����oN�e�������h��k���/>>K��f!5*��k�`�PI������Ơ���u��C7=]o�O�C�l �B���^���lr�I%N��W,.k��kPRg�
����^O��㝈�3>X���q^�B�Ux�͘����U�>
�����h�k�z�k�Œ���S{q/�,�����a������:�1�AH�b�S���-��W�erNghNWn~ј����;�X�.;�r֐,gIr���O�Z+#`��!Vn�8م�fg2���������%e%���|oƋ;/��R&�X,�=E���r������$��<���s��{�'h�2g}<�����6 $��Oj>���:�������׆[��1�~�� �$��,ʪ���[���<���ݚR��:9�����m�'��r�8Y�HJ�ƾ�\n�q\�8�#k�Qh�֍D�.�BN�rX=E�$~��-]{�L:à8J���Nk�Ew�ID�%�0v��g��;�����J�lw!�M��#��� :�s���E�;�g�mW�5��뭜�|��kG��+s)H�+���<��:����*��p׋ڤ���h���%9�:?6A�Y�|!v��}��v��^=�����7��:@9h�Z#_��<%��Qg%��(�ԭ�*j�sP��o���o.��'8��'̷ߘ��0��e������-����V5���> *166��ge}�#,,�́���<y�9��z>�IȚ�m�9F  �J>_�M�TC�3�+��a�;[H�s@���7��e��T�r�P����/�����rU"�h^� ƭB�ؽ��簀����S�ɝ>w6�0���:�K*\o�e���>����2�	%�G0��ҍ�?t���Q&�N}����1L��Ŧ����T���ᆚ�L>����^?���2��_j��i�߫N>���/�N�x�uv�V�NA�g+��{]��� ����u7��3���t���I��&L���.��������`��/m-�a�%=�큡�8o�뵻�a���㑬�@י��&iiIh�^X���OVso44�%��M��2F^ |zrlp��"=���pJ
v[��N�t�0j��M��f�0����� �W�Ltv[�!���).�ɚ�n�	۴*��[�+"��v�1SI�L��ص�ʯ��&8-�S$���7_�6�t��Ӏ���Wy5^��\�2���*v7�/���?�h8��������byw���I�΂��v�	ֶ|̈́j���MYgb{u����U�~!%)��Y��t�y���� ��5�Ny�'݃qq���z�5P�4�4=�5	 SBئ��/��aEWF�_��i߂2tm���:7�sff�]�,|�����-cšt	X8~�����Cw?���QF8U����L��J��$����O:�-��e��4疤��У(�J���1�df��	�v0N}�,�VWp�|�ݢoi�@�iQ�8]F$��S�b���<����]�����dU)����1|�1ǤJdd�I��aУ�����M"��C��L�V��{�e�D����ƶ�Ł?�D�u# �#�w���Hۦ�û/��$��Ia�h��6}qN���+i���A���� ;=mqQC��+��~�Q.�S:��W���­n���%�1םlp�����C������q���" �齖81���/�(��Ay� �}��w�G�!QQK3��f�bͩo#��;��n�W�5na�<��l�>�{aռ^��8܌�'nXO����cN�/��w� י�h�)hc����$��Q�i�G.�1G�j����KS�]ryE���ۋ��m{h������+Jd���h���C�i}�G�ZR\��+�ܙ�+���r�9���r#0YC!&]��W˰?�K�]L8V#h4Cjˎ78��N���3�7�F��7�&M`�D�3x�&K5����O\�B|ef�|��qS{�5ccIeݙ;o�gbV�o��bŜ�3�!տ٩u�	��P'��y�ߪ���XO��;����
�<���Ӱ@��l��}����ON蠒Y9!"����4���r}���B��{%�<�Dֹ	q�����5�l����m��i�?}b�=u���ϡ16f[�艔7���1ۙ�ƙ�޺3�n�71}c��ڙp��* d3�{A�]N�w$�t��!~���=H�t@ۨx�����`Wr���{��z��8��8]����?����ȷ1s�
��V�VFk�[0<T�0I��*g�z+r2 ��I����%��4#�8N��\R�����K�Z��/D!�;f�$M�\P!!a�ЄT>�Ȃ���{Zg������z�m��ڌOO��-ʓ��*Ch�����=�[��Z�HN�'0�d1?k���F��;ߍ�ݕ�bv��SPF:�af���oYZ!@ȊJ�Y%Fά�v� ͤ�n����x���_< �kĵ�\���/�9V�Ky��o�z�����wOS������o��3�Vi�������'��������G c֬�+�sqW�к�D5��n�e݇��o9�7���\9:�������$���<�Nh��o���C�^���� o�x�݌r�Y���ַ�g��K;���s�,&i��i��L�D��=3�w�F;�ϔ]O[���>�!<f\/��'ػ���o͑tA�-��h�6��x�/[>�wvA}���ge�p'K$T)�C�,>oJY�K#a8g���h���e:o����]�����Ŕ��JT���8����H: �ڞV~ϛ�;p���n x���&G�����������"1}���Nv��Q�����kyt�4S��<c']���5nn�;�W/[df�����3��R��^���+��� �0�	(��E,qR��ٝ�pz�Ү�
pX;l��&�(s SG��� &�=�;��P�9�7�+�8���ªV_�VP0�2}ǙR��8����H����[E\*�l�l���_n�פ�A7%���㫞����g_}�]��1~�����	�� ��}�Xb!�&����NDo�����7��X����;�~��A����"^�mk��e�?�X�碌����98�By�?�b�g��1��s��v�6��a��-^rh ��>!�RF�"@�Tj\���. 6.ކ��S��a���i�@��DV���~��g/��n$��<P��y�q����}p�J�K��u�AE���VX(��"΂~1��1�yf�>HDAx���l�$Df�,*�%*Jk"��e2G���3�	5���1�����*��e�x�=�׻hD�74�ԇ�<�C��2�B�ԋ�@�]�M볁�4�In;q���t[w2 4@�(eF���>=@9^�,_�{��M߃�O���y�Ω2�C��W�s���5��~��
ķ>]�I!��	��a��D��V�t�R]%�Wh�`�'�AkD�l�#c⹻e�\NS��2�+Q�M�
wL�lB�γJX��Һ�[�)�@��R�Z�>�L]�U\F�fF(_��D�m��5�s�:u�qq�)l�5�9AR��#o�A�����tϸ������0�Ah���<̡��T�$B����/�%�煡��������'[ܰL	����	\Jy	��n+Q\�?��g]ol��[�Y)J�\�hF��d���	�g�mD'�G�{xٝ���vN��_J2�����\|0ש��ԓ�w�`ΐ��㞧�%�1�|�jm����@�_Ƹ �[��C$E{�=�57^//�R|6r�a2�ϋ+-
� ��F��	-���i����P�b;/��W��6��㹔#���:Ƀp9 ͒����0Fmf�ώ"􆈐1�̡�[n���e�5Q%��
��9�=x�e�.���IA��Ǳ܆uwK膣Ezd��a�w�l�={��YӍ��>L2�z�xl�|D��i����%,��kv�QG��t���n��J)����`��l�n8e�Ϻk�'|��ځG��|G^[Ա���L���އ��x���m4��(r�xU$��O��A���8'�ثD����k��?@҂Y_h<�!4�Ɨ]�/V�+g���>�4J���J�}�x�VPF8c���±zA��̋M��g�|d��d����~FiL��cA�j��%�@>c:�+��Fk�0{�,.�ֶi^� �(y����>p�sSx�=;;���yѿ3[+X�qo�Hql^�[o�gvGN�uM�/��f}���Is��F�*-S˟F�}�H�k{�}a��`"�d��OT����3��A�hy	O�;g��ZlS@�D��Q���;%bo�6ƞ��hg#E�U_��F�A�tH7�)
H)�).H��(]��t�t#���� -Ͳ�t.������;�2���>���|��y^N�:>�?�+�mi�|��eA>TߠT��~0??�̟�o�~�	��~�>�������d�;]���W=���w����Vɳ�zKs�_�F�,~"`S��u�kRA����4�5>���%	��_���~b9�+0_u4�:8�h!w\������c�졏��'�e]L?K\��5���vN[<�u��H���ʍ���{�gU�L���b�PD�#V�	�9j1�F�|���qv̛���u˪��Of��fQ-Q3�)����QJ�T�5�t�lR�]D�`qÝ_�Vۗ�O���,n��X4���u���	h���O&	:e����JZ�$al�}g�H�#iQ��@��3I�����F���&�7�lFq�	g�5j�Ky��1�&�z"����
Oz��^(x8�%� ����+�M���%lm�}��N��w�ҍtw����r�C�/�q��̖��Gs���`G�k�u�!)�V�z4�����j�%��+�д��f��/���j��K��w�����nj�l���ߴ�����+�W�x���2/�p�r|�=a�b��'��g�����*������d����o*�d���x����f�ec�
`0F@���]�_cZ�i����=<���$�	��>l+}����7}�u�퓍�U��(�.�OO؞����0ER/�`�0^G��,���Oz=!o�X1��r�z�g	��ڊ\�����*k��K/K���/�g8�����{�./O��O��`n�&M�ۃ�+W��ʬI����B�0� n��+�
ד�F���ʌ	*�~��3O�/�G�J	�1X�-�����A��nͼc�zXF�i�7�C2�/e�6���N���#�6ǸfS&�_9K2*���9��PU� ����pA	��oO��
�6wB7��xK���3�TjĊ#��0y�H#*�[����.�V��v]�x�>r�Ű�w,L%���G������*wh�QĜ��i`vl�ߛg�k$�=	o{�֝��eo&=�.�g&�Ұ�l�lﷵ(/���4��+O�0l�Rݥ��`��$S�V�<�LtҁtWJ!�f�9�o�������bf�u�&��kjK뉢�̡L/Z���0;��L��������+שmwZ�2���4xl�;)�8{e�'j ��ۣ�M���:=�.T�Ѐ��H��0�.��������1ܗ�L��ó�?�/�F;׍��J�iᗕ͠�M�
��-��J��	 � ��1J����ܢ��NJ%Ծ��4M��`!�>�>⨞u~қ�)��S���V@tt����:��'%%7촋F׷�F���}Q~@W��٠�lXǏ�A�Ȝ��j.�Q�'��y�����'%%a`t)���	RNz�1���?n�>��*v��b>��� �/��1������K���l���p}���r�MҪ��؛�-{�9�R��S��﬎��Xzׯ_�5]rH$r\��֜Q���v"--��2�Z���}P+n�&�=�U�bV�}ʫ��yN�7��zh3�O
�Z.�:��̗�Gmٔ=�D��o\c����3�4���18��;����o��?�`��>�>���B�s�(�]����ǃHܦN]$��R���	�!Ѓ�RD�G�/q5k��z�$�L��zj�3�5�t�%**ՠ�}�ֱ��8"˞�c�Joo���`8]r�E�� �v�e,t3B�sn���\Џfu��ҨX��9�0��>=q�Oc��7��/�(��j?r�������I`� 3L
��Sϱzܵ�>n�
 ���'ω~h�9K����$��yм���U�e^s	����,�b��u�+�G�Rn�<A�m+�F�V�3R2�9D�:��̇�������桁�\�G=#��R^jglKn���w`խ���+����w�^[y|�(�SU����������6�����+���er����7�.�&�m4�wu�5M�^� v�I�((��}�ޣ\���=n�)���-�L#�h�dۋG?\����4�4O������
�	�*s|Q����9��J��~:��^��ߟ�Z���$G�G��]��Z�.3�E�_`����O���,�PN$=��,��4P��y��u�K�~�;(�|m2��|!qT�!_	�gy{7�� �^:�1{`�J7!:��'��\T�zA��İ�����/�N��*�j!�&��xG栗RP��=�=#�aΣ�W	J�۫NT���Y�z���hr'/It�J���T�{����u��@j|�;��N��b��S��?�ң�?8��f0g��t���%�d�s�$*����ћU���B���٭��?����5���uӼ��ʀ��r���W�Ύ#9&��ݗ��]�ß(Te���^���qG�E`T�Ys�Ik�Pgp���B�L�rt`z�g�h༖������ך����3Skf�ד+�g�M:rHZ���l��'sxyw�5��< �d�&br��/���x�߈S��Ⱥ��Q�g����JK��CV�V��)��e�u*�҅�02�a�[0����c�n��hz�|(��@�9�/��^X0=��%���x������.a����m��UQ��&0��?�[�yy��� ����	fMϵ�ټ��<ݩ����]8�Z����������fD#���I؁�ɺ���8+nӆ7�X����α z����D��yL����L���ͪ��S���� ��������(2NAQ��#_,���Z1=e%��;�QPS�ۯo�@֤^���Sֆ�&l�(�+�O����hf�W1t�J�������SW��-�]����_4Н�a������"��/�;;Y�C��4��0CTf�-���-%��L����ϊ�`�.���I���G򀿖N�>V��gK&����4mx�x�j���.��5p�J�^�)帯�A�1Pm�?�	��QjP�֫���ο1�4x���|�?�d��&�V��cA�M�IR������)����f��ͫWM.	/)�<znӭH�uuuj��[x�����OA�WC���˽_ ���lf�bIX<�_~��
��������t�)�b�T7��ñG>�{~s7}�1��b����W(�+˿["8Iq��h���	j����n�����@M�/��c��9�*"}�/��jS~P�8�{���r��o��
�K��^���ٞv�K�Z�׎���(�����	$�ڟ��6�_$������	8��TZ�d��z,6Y蘿��	�#������kX�BЗ@��g����=_�0˩�p�KJB"y�/����D| �f���u�sj���t��s)�7��U(:�֪֡f��ww���M��l��?���U�>��R=�~x�zG��W��~�d�e�ե���s���6���y��p���d\=QB�_B�d#�L��3��]2m&�i;~��2Iqѭ˴�D$$p�����i�&UC3���.6��Z�!�હ���+�v~�X��o���O�N �P��K����$��&S�ne��25/�v�$�q��az��ʾ�d8eU /�iT<��bmt�%H�M�����Ә�p%oP���k�|�8���m����qS�4H��^��bLb�2��Tط�nX����?�u���z\�Pe��U�<�Ү}��DZ���C?v�*!��4̢t~j���E��O�?���2tG�F?f�T�avW&��\%��B6q_W�L_���B�ޢ���ۈo�vj��X���2
�u�x��g��ҵ�ǷL�C�sS������q����8��|	.�mX���}�D�u��Y���mʃ�K��[2�d��>���;z�J�����?7;�%�htf��y�j%����=Ce����E�0ڳ�clek|��J��b#�m��ҹ�����A��]��C�[��sD7��j��;�)H��^oMb�����Z��w�U�x��Ȅ�fP@`1;�L}��mp7�A�����:Qx�9~��i�8tvLH�˔���t�P�� ��)���Y�㍝�S��ț�N"Moӛw���ulm�"��>k�x��AgOlpr����I�;��u}�w!\*c���.�(~SV)1�����������t�O�V�a���`��8�����,9�+����z����sA"}K�n<pd}?���Rz��!�&�t���b������So�ĢP~���ë>$c��M[�R����=���k��'���G�`�bg�����\i����B���Dڂyn�R��2K�Ϗ��Vwn�����2b�a+�`uˮ�o�$H��������ӾR�ܱ�D���$��%��G<�R�fj-���X�-�RJm�H��{��8��XI�$qj)9�A�/�~+�(y\2Be��=��@�5O��J���/�9$wq`�{�-����^���0�vzv6�{{��+�I�[�rE	�y�s�Z�G7�z�$�[CXgwQ)��C�b���B�����P�u�%Fq�Ge����)��usV|�eCRB-n
Ov�ަ#���y'O�}��	]v����%a;CD>�S��[��3�RN�!	$�:����XR5�\vI\�t�/��*��A]��<��}��Ŭݞe@���_Cg��l����]m���Z��YA2�9:hZ�$g��R�47��5��(.�@�XtJ
~��m.���s龺ݹ��$5���\J�1�Ҽ#`����n�K�V�Mq"�X<�V�9�8��n��/D��6r?��J��gV8޶�V�T�z������"[lf,�'G�����U�����Խ%jo0k��@��hM�"��Na3��s�o�x����a���1�&�vv.05;{�	o��q�r���Xս�7aByF�\�W/�Z��vv�|�C�(K��ڸGts����Z����0�c����as�}]0g����	�{�@��KM��l���lr�1rx����6��e�r�JL.Ԯ!�PBϩUpxTi�?����_�*B1��_"^���~�2��fO� ��h�~�.�����8�쵺=���V�K�6Oe�%�e���(I�#���t�t�!)��"@W��oN�6��Do�/��J��o�B�,��W��gBKʘ2�Y��<O���/�̓�����Ѭ��� �_[�k|ef��;�o� E��]o��2r���^����y�߁z����kh�~W�}�LwG�݋ɞ�M����^D�9�M����k�_����~Ҏ#+w6�(1ѿ�]����+��d���Q��L�X<��Um�/
w[4(��CR�t�@L���f�.|o��VO�A�6K�IG%\���Df������ck��)_*����4�{���k?���j��NrЏC�%�o:��(�xH}��fX�:��I]�Z���sN޾�:�����������o�LDtW���r���;e控\�wk��X���l���w��l�����$-����v�;�J�BW��!4���H�S5��s~/���vg-(�^eċF@I�6�NfȞ�l�>�>�kd��9����z)�������JEOO�{C�y��ig�6¼���rglt�I�ުZ��n]E:\�3�<�j���6�s��W���I��M�qK�"����e90����W����c\LD��g}���H��=�`O���o����)f���96v�S�ۅ��%�>$��-~�?-5��1��E�$��ޡ�&�8��9���ou2<��U�lݔiH�����cz�=	�K���c���'��d'E�F+�WM7�0*iկt�I�[T3C*��~�	p1���s��v'�_�|�u�:�Y���u�B��T��T�k}���Q�O��:s�����
r��w��)�wf"�^E!�C|�&��B�J� .��.�}\X���tB1�៙��f��W�L��U���*wPki=*�3���q�i��)�rN`m"��3�$^3��X�d�����o��n���<�����x��,h>t���� MT`�W���0%gp|���Ԓ!F��}�ao� Z�^!�Zx�p��-�fM�U�E#(�����˦`����&)��沌�K4�h�,{~d�ϫGߍ������K�m�^NVA3>����D-����Sծ����'y���������([��88h3�h��`@lH�o�k�P�шG�@U�y���k2���U�D �lȓл3��,�!���������ZR�E�-z1�_NT��؎��De���,5�$�����z:�g�z8����į����G��j�'�tuu#�8B��p4G�f1m��ނb5oW���s:Sc�Fm�|�D��эT��^N�Laʣ��H�x��є7�u>eh`�j4� !T񋋨ܢ��%�������C_���)���jC�+�J��z��bk���H$>�wû�➸,Z�x���K.�lV��D�� j���W�BE�6~�e���Ncͧ���Ks8xj"�KՈ�w52�
x�&6���yl�P���ow^�I%X�#�h��ݨ��W�B?�͘m���pOPH��+6�����L�7��[n�Td��)��C�௦���3:���/}�Ĥ�^��!���,7�譀�E�e�#g�̯I���.���S��6���5�c�<K$��0mI9#u�����?C�ȶ�٣�B� �m�����\���Ob�wIȊ���L��+(�dw߱���1���ߝ������0�r�n/{N`��s��r�~afV!E|%0P�L���+�o+$���I}4�mv��9\�J5~jB�vk��q��;�?X���ᩒ9/�ð~H�7�((�6�6w�����W�'�s��	���Iț�?�7�B�T��8���o	}7yҏ�_�qR3 ފ��poC����sΤ1��E�x���8%d��T�Q�[B߈��tW��8e���	]����iS�I�� �Sv��U�Y�$��5��0?T�
I����^��UA��^B���K��׸��R��c��K46��Kw��4��`�+�
��'����튍�8���t��N�4Se{�0���&�^����8�ק\��EBe��0�����,��!����
Ǝ��\B!���&�!�X�4�zw���>�|��3ڬJ��H�-s���g�/���=��}Z1������|Qbb�]�k����ڡ��|���N#��+wr?�
�i�����`��$x@��!�mEg���1�,Q��f�1�dswY��.�an�'\�;b�,Sh�dG5FPL��v���0 ��H	WVV�Z���[5�p�L,L���Q\�'=YIH�����wk�kD�n�<����L�j���C�.ںl���ġ�UvP�Xp�s ˩���qB?��� Ōf���`����6��^S�oꪒ������h�P�\�鿼���;���f��
�s�����}���y�PyѪ�.y�������N�i�+�Mxk��w�<߯j3C<]<��O�p� ���A=��<��ތ12�(���W!����h<d��Ӽ��.�̭�g�?�Hgc҂�ؙ����d垝��K�sʬ����)�rf6!M?/��3|�g�w<쩤�"1Y�̨�!�������@P�ʱ�$��}das�2���Wפ�w�M?E˿ҿ�a:�4�ů�/��L,�����G+�-7�@/�~2�ؒS>�Ǧ������;c�=��Lݓ�. ��"�ܦh�J�A�d}-͔�ʔ�k�yF_�l��DRٺ�G�3������1#vc�� �8��^�6=��8m�.A
�4oY9-����q�_���l~��:���k�� �1�_i�|�/.���"��Ռ�?�c�}���p������_O�x����!�6K��5wqQ�5��<���/)���2$%L+��������ء���L���RM�޸��g)����?>zA����������r��m��KL�c�&<��s)`݆���.��r���6mI	5i�D��4�_���o��x	�bO��ʯ�av��T �	?`�c�?�$K����KD�ۇ�a=���yRm9�7�i,���n��oO7�j��Y-gH�o)K��D&�q����#P�f�?��L���Q����C���}�7��$\��ր�ш���S���,���J��oʸ$�g3�ŏeԌ���}��Ny�����/h�HiU]ޥ�W�Na���`պ��o�3�2���]l�/�6"���V��D����o��z�����Ï'��<�)4l�
n��{H���Ҳ�+nm�^I�?����<>R���}N �
xǧ]e{'в�U�z��ן)M���+kt*�
#�5����� I# *��:�L�m��#��(����)jH��z܆R12�D�-��y Udx�cI�� ���6ZA7�s��\����/�!�p�=Mf+�9h0[2��-��u8�y �AbT>G����Fx!(㾡ߠ�`#`��[�)1�p���̦���-o�ct§`O��YT`��GTM��C棞|�򋷵�0pQ*`t&�65�T�w��I����9��B�����I
=U�;6x3O)�v�����cD&���כ�ұ���5���r�z��l7��s/3�r�J��0�<������������"TC�"'�p6�f����(z�q��m�N�;�-���/�a��W�����I��t�pf�HQh'��*�2��%���"f���;���������q��J�	`,WJG#����RO"s4���"�/H��Yl���8�������("�KbY�{�ۛi����a�����]�|ӆ���ndd��~'�!��D�ˌU[��ޔ�8���8��Z64d]���fH��S�D�����J1P$�`u��5��H ��F" RS9���IQ��.�Q�砬�2�:B��-�ȃ�s���ܾ�K���T��x���+Aw6᲍ݭΘ�!@Ʒ����"Z�}�rM�@�]Z��Y2h���٩A���O<���!�S�d�Ƕ4y��##8g���<j~�f7S������C���5X�Ϟ�Ȳ�ʝ�g ��&w�����N�5�X���lܯv��X0��M��-9�}yԫ���&ɦ���T&Џ���x�î6�	��hۼz��\��T�#"�xҭK���M�gI��p�Ͽ��9��Q++��B!�"��M���|�b��h�*O�J��f��ު}}u��Y�@�M�!##P��]�b@�um���O���DT�FKG��*�VH��|�L�=�نm),:�5l�E.�L�7!��v�������vM�ߩ�c�S@ޜ���-,:�MQ"B$���@�jo����DG� C}��Ϟ=s��.Y�t�ś��ݑ���e��;�O�x~���K��y�x��~"�30�k�e�[�$���(�_�--M*�pH�����e烏7 6�����,v9G\�{H
tJJ�D`�"�W�ؙ����Եy$�;�&=���B���A1���CNa[��"�s��u��}l��2�,�C߻<ȁ�����|�s�>���B�_Bߛ��W�BNr{��Kn��v�zV��`�@�$Ӟ|���90�j�&��F9x�[�D
'I�S��|RS~��N�;p�>kǳ���fj�����lѧy��vl���
��q�G��|m����ǂ��̬%�t0o���۸P�<������p���MyQ�p�^��V��M����pKy��'M1��A��������صq�٘���Om�ޚ���?��b%K��ӆ�U+�d��O���Y������Ŧb3D��L�����FT�3W)���̮o<��c�
���|�K�lh�`����FF���|��26��L˛���'�$P���CRrZ���5�<$��l����^
� >j������
�@FMV�������f##����oU}�?c��˪w��о�A�s鐮4�����BI����F@+��T�z	1Q�>�U��o���z֒����Q߬�iC6�m��(NvT�� ��U����ɴ9�����H�k��W�I��^���8,��m��}X0��F�MNB� &=-�����d�󬏪�yϛ�5����������
NQg��ɰja�`���:��f��,f�̀!�Q�-�q)�'fJ�4o��	�-[���Yb�O �T}o/ i���Ч2���ÞH ��^�o�f5��� ^B̩dҧ�w�^Ǯ��������
��`���!B_B����.x?_��Ĺ��_�'i�_�����Ʃ
v?��]����������q�o3|H��P��2$�|��[kl�iQ9�,�������&J�@U��w̌�Nn��un�-����[<�����x��^'8�����I6��"��V������`6$��0�������G����U��3Q��x&�}B����ǂ�� JbXV=)�i�/F�[��8��7#�cF[e�==@iՁ����u�/z��M�6�PH C�C��p��~{�g�n�`C*�s���$5����͕�`��T�M�wm��Kv���)B��٦ |�$ގŮ�"�S��N&[�:�?_驺g���H��
rssf�YL�ͧhYA&{��+aǊ7�������e��-? ���M!����"�r{f��A�������r�	�"���6CZW�o�7f�!�Owf�)/hz�gQ(�r��{;	@����}Q��8�)-+C �5�*��z��iK E~>(8R�r��3�'����|��M�6�T@���1m2���R��.Z^"*����N��IT���y
*e�\����K2�u������/�4�*�����j|�}M��n��6��Y1T
ȯFR��	~y�a�x+��裢/��biUl?�E��������)�uo[�����Gm"�˟M��O,VV��;z�؏�b?���&�l��^�'
�'{\>�6�f�H8��&�}������F$-�,�	ȏ�����]�S��;�Q�,�.����� bLj�&�۽���L���1"���T���2��0���.���TS���s
��;8���sC��4G]���L�[����ҭ%?�խ�ݩ�h`(
��w>�f��	��TÓ��[ǭ���'{��8��dP�55��C���<���� ����U�Rs¬�ͻ��/FEBI�r�_����P�~�H[#�*&�y��^�{H��6 ~{�{�%�s:V
xN.���߭�X-g�醍N��iܪ�g�T㕁�;��h��xG ��[�UW.}H���߁ر�IϳۢӾ�������ls���V������"�Ņ;&�+OƏZ�o�I/��<�ř��G�r�j)�S�GP~��d��~f֋߂�~c� x|~yy?=�ݭ���-,(�����	�3�2���KVD���.J�����Ӓ����V�l�;�H��1�Y"
+��Yj��OX���uu�B���b�t�����!ֿ[/��Ҟղ=�'�3�>9�0�$�pf�P~_u�T�����񛚇c�N����9��<mQ}��1E�&�V���uboM��gk�-*kg����MQ�� x\sPfq%��ۦg�,L`f�V$g�&�ܴ$��cg�KcQ辪ݒ�C�����}��<�0M�@����v�F�-W&��sc�A�M�����vo���4�@�S"���ʝ�����۟Ar k�2�`?%��.����Y\f�mDLazd~�َ�w��hF���F<�]�)�O͡������Q�Qp�Ic��wnY�w�W#���gC~ȟb$������4݄�0=T2��f��:gb]�h���_h�/yJx�1}�ʹV�(\��7i׾���ѥ����/-/))iW1[*)�4:���Sĵ��ig���N⓸����������}��G&"�+s(Sq��:���`�����]5q,֥���B�i+ݟ�~���)�߮�M"�koW�t��dsT�KF �	�lc���w�"A�����ˏ1��}�Ɇ��z�-��h�!�Ϗ�"���y����A��H�ڏ&gC������F�v�n/�5��W�69.�ǯ�oQY�.B�[q\?�P+d6�)굿����-�;���v��bs1���'X��-�<�,v�������)�g�Y�H�Q����4�B����蝧���6=��O���}��?�O~�a2�WPX&��'C^�S�b����VU�ʏ�+�"yg������2�K�Yg�z
:aP�"����_m?ا2b�r�'(�R���*�f�r'�f>[HPP�X�Ր�����qR�������r��J�Np  �O�#�B2�AQC�S�����P�ϖ[��s��URҜ&x>���}b�gsl�'r�7�y�Ec�IM4*wt����p���kE�G����"y��\B۹60?XK'��t�H�����ة��B,"���	�^�dcB۴U�Gh�+Iw����,������g���l4���a���MQU��-���Q��f�_�~�)�0�䵴�]<؆�g�ZRߎPK��Þf�4u ���Y�\z t��(�g����c	�91e;�x8j����ڭ���.?`[\�(=J��rRy ��q�^j��F*Δ�@J$��rՙ�+�
�Z��ׂ(ORH���-q��+��w:�l�D���D�~���층���0�`]�J�i�VG6�Y�Q�}#[ku��FR���wT|yy�e���A���=>��=tc���[-����~����˦�"5�����G����T��)ξ~~�W�*�ff����aJ+6�����:%�:%_?��z����=oiKPT�M�����o��XN�˓�A5<�u�Jj����E���,''7���}��}f!y��Ԟ���K�'�O23��1��?\�/���Zj��kp�ڥ�b��r�PJ/���p���ۗ,����#	=�f��d����^���!�����-S��j���O�@����>����s9��%�kF֚�f�L����[�d�PlE(���v=t���B� �����i{��s�0�zEG<郮V�Ov�#�Z�6%�פ�7Cm���1��
�ϩ�?0��/3��T�n��=U��>y'-d׼Y�*Ruj*�A������cM�����b�WɈ�( �$T56q��&'�/d���c
W�uzcO��Ч�K���Upb�ׯL�ϹȠw,,���\�5֐Xܠh�&Ƨg�В#�77�D&�9����_ۯ�
���1�{^���e�T�B�o,C���빼�#]Mc����D��"EϮ�~�6�vXPN��
� �����OGp<�����*X���(�r�\��,��¨�s_�����R����k땯���ŗ�KKK�����U��V�����C�M�66�w�?�u���z<�e�{�-b�w��G�uuq����匎��g+Lͼg7��I���A�%�1��	b����2q^n���T.��R3���K�-ǎ�����L]ZZ��:��?���=$@s��!�pe��kcG�]D?���1���6��9�˝��������I����ЫgILc�h=�A�>����1n� ���h˵g_qZf���/��F<��M�>*Z��eq�3)`ڝ�M�@���ƹ����:���;��|?���[R��Å�e�����,x-N���'��k��Q�M;�i�gҧ�>a�HABB�����]�Ԕ�뗠�guC)J�;?�X	G���/ܜ�<��d�+��:Y�R�z�6����p��������4E:%\��x��  f��s�gk��;z� C�*#.��/�]Er1kBi��!�o�&��[���ʅ�I�k�Z�x�̃a~��	���a�2�d�,�Mj�b7�����d�@��O	�����e �F"���V1\��=N��o�bz�E�/�J��{��D$ͧ;ס�/�Q*ϞˋF:î�n�.�b��c���*�������/΋�D�T�%.�uי�[^� \�w�4�q�+/�i���`f��/�49��Na�D�!5��b�&<���,�mHe~m)̀��ڿ�½3����'�wƖe {e˅��ݹ�G�FMԀ�{�7��	ikV��*G���j���b���SE8��e�>�A�uK��5�4Z>m{HϠ ��4�Wċ�5����	9�J�`+�����P��B=�0867���N�[�P�^�
vo��3f�L�5]%i��)���m>^HT4��p����47w��@��C5^?P�^��ş㶢:|c�3�O'M²[?-���g��o}}}	ZE��9��NP�dSII	�Q:�ysl�p�h�H����$����BM05(J�FT�319L�"��Q��>^U:���	N֐q�0e��ƚ�6�E��K/�:�a�xF��@R���3̝��a�X���H��'����L�s�=��⦸IE51)�.��p���ƷC����<��q�E+�eJ+���p�}y i��=�M�.��uN�3�9�r9?�?��rT��SЩU�"Z頳(;�F�*\�j��<߸�=���q�|w~�G~s��8��5ݿs��1Y��㞄dǑ]�6i8M�E�?��2��ňw��v�4�9�S�9�>���)H j+�"�GMO��Y�0�`�h����~�^;ȏ�ZWz��M�Ǿ�Lj�^��(뾤��Ѭ��*G��	�L����m��#t������+Td���Y�Y8�8V��ER�`lQI�4�g�7��!6C�f�o�j@�Xח���
���W��b��XϓO�`G0�b�t�a��e�.DMٳAĜr�+++�'�8�
����O�%�h N�:�F�?IO�%OP�b��j�
ʪ�x?;*���I�j��� ��W�D2���Kdzy4���!�)��IŬq���1�r���� kq���,f�љp���u{۟)Y>����oB����{B��^��[ �A�w��v==�o���ill��*���H-�W�@���8[� �]���F&�r������#�2�+<�S��_�4�Fv���4`�6�t
�j!��9���#�{��_��+a��.��X.�~ᴸ*�������3ҩ�e�pi��=�,�x��B��ژA�ej��2N�_i�(��R��M��1P��㸉��r�=�r��� ���ݮgn�M�YJY�6*d�mK��[��'���;Y��4?�����<��LK:�s@g��il('?�*.¦���6���7kw�BJ��Y�����݆͔gw44�M�0�&R?55�>���p��6�dQP=��e�g��%�&E&7WCX__���O�%UU��L�΍/�FZ�*���?�����W�@�g��t0�ǭϷG�x"��l��.+ߘ��G�ES��(�;ȝ^<����LO���'*�~�Y[����%x<kb���ic�՗��c�fy:dmL�.��)��x�b͕�߿���o��:~�B�z��3��%�_0�'(D��)�
6b<u�Zm�)��,ە��nk[/�9�c�[4��E��i��JOX������s���5���ڤ�4�Q��� � |X\�no!1�s^�C�w���'-�C��k�>�l������pձ��m��R��~b`<����Xud͵��W�i0���L��5Ng����5�E=?�h�V�5�ޱC��W/�,�~7��$�U~\ss>��$QO�|1*�x��2�JD�J2����]�XW���}�͔�'dz���Q��g�Ⓠ���]�fл+JyK���N�&�c�b{?s��\L����w�s�^H��I���p�T��������V�~(��խM���s�4����m�`�y-���P������^#�[/��m �%矁�=2l�lp���'-y�x���w���]/�Fm��w�% ,N�;�Ⱥ�ե�'>����>�=�z���߶�xk]������s�����(K#�H�Ji/uj&u��]�P�dEW0&�ߙ��B�pz'��|7���?��U%Z!:��Ѭ*q�:ؽ/J03�_"��
Z��Y�2��<iA��)&��ڛ��iO����o�,R�q�t�cv"X'��ɴP�py�����I{��g5U/�elT�2<�b2��������0��ppC���v�t4+«���LsG�FU�.�A��q��*kj>���M����3 �F��#ej/TU�[=���z��e�N%���G������RS�DZ g�7a��{!|��p�R�޺�	� ƽi����1���}{[��&�$���pJ��B���C2FG�M�F\��.<��6�rlR�P����\ �����6-�~��VQ�'��O��&�0�,R��Y$�.� ��Q�����	|Y�Ђ5/�x�YB#,���q�MD��Gإ5�t�+}���P���i�������ƕ�uz ��q)
�o{���5�c��qf�n�TgQ�4k+� ��׍��Я"�w�ъ�[�iŤmt��ۅ��B����	tQ�y��!��g� N�U��EY׈� 4qȩ�_�Q��;�ׯ��y���'��ǫ�X�Ť�]�p�;��K&I�;N��ޮ��ωK��o߅�H̶�9��ɛ�F���D�oW]^�O��TEj��,C�?	֌��z�t{��F^6@u��b�jH�H�-���~�pK
����
=6&r{,&�i�X��tꦌ��5l[�,�U�9������v�, �l��K�B;ś1�u�l���MgVzU��W�"x�o����Svе��,�����ͽ�{��&p����2U�C���XO��A�������چQBR��Q��NA�Aah��SJ�N钆A:��.)��n���������pf]�>c���M�5�*Ua�~�p��2#�wJ6��1��,:1�$����
����j�i�}ϣ�A{�n8!��x�J�ۿC���)�CTXXX�v(QktD����腩l~�}�����d�d�Q�:���U
��?���\��e��74��kqc���DFm��a�~��A��",�
P�b�p����/,��k
��\��ٮ- ˲��|�.���2��sV9��|�(�Ӌz�nd�Z�ۤO�c#}/��'���^������f"m���hd��V��s C�}C���sD��)�$<�=�>l�7��(�1~�8~�ȝ��\���ƀˠ�ͫ?q������S�z� tt�!B��2���&Y��Z�������z������G�#F�E,�3n�xe)�w�Yۄ �)��]�B
(LC�����L����I��e��F�+�'�xiv����OmZ��C]����`�v�G�\_v��a�y)��{~O��H�	F^��KS���/]G�l3ª M��%�^���ῥ�n_�Ev���pw�?T���N1�2HǨWR�gv��z�A2��W�bM�$j�~����n��n>�b]�`�a@~��`o���l^ e|a�?D ��Y��1�`��N�8�n� �o��/1v>�Q��.� �>�_�?D�rQ��H;�cK���i*x��G�C�O��7$����j�����6
��(?��\ ���bo�&+"� lD�G��\���֣f��;Q�N��v+H��ijc���$��K��S<;D�>V�����R^�Ƥ ���5��(�p	�����(��ܕS����,6}k������?1%�9��j:�t`2��h���!×��:vuۚ�E��Nc^#q��P����Q#����;��B�_}cn.B��V}��A�
�%�77�l��Ǒ��|��.߾���"����������>-�ã:}�#��x����HrWG�B322�N@	�^�H�\.9��\I�^%~	�0-T�(l����d����8�?�KlőD���[��d��ϼ� ��������Y]�}6���O���D��u3i�`_�j�vM�?)�HHͣ5ƿ�,+32(���3p_��ӊ��V�O�%�+����ܡ������ I^	�(@+�%�;K�K#~�}����9Gʧ\�b5������-eaX��^J�wP���9�鮀=ےW����S��~q�/���킼�CAV�^w$����Mwg\�:��g����'�i�]}��#?m�s��']�N^:Bۘ�5.�w=�7�� U��X�������"|�QbW�.�׼���wp��4<<�1����I���&�
?7�"����U"�U�t��́�p|bj:T��A<)Sx�Y��c/�4��Y�.]屫Ӹ㵐��G�X�s�]5��'�`����wz��},��n�|)#D#��J�%�ġ�X���������>R�W�N�Y^!ۭ�U�b�z��H*��s}�O��i��[^����k����s2r����p���*U6d�����g��ݎ�_�W;6̴,�J��h�zNj��y���&>����`�u���!wiZ����f�߳1�i��اy�\��4����))K�����:	�K���kR.�@�>�����js���K>����x�JD�"���R�����M"����!u!�����^� #�����l��2���Kp�Q��mX��;)��xn{:�����Z�%W�B�	<�����}��?�1<O뚂�bk�&p�@���/��eCJ#�]*��<�A��p�P���Р�!��ɰŕY��M*K0�W"��7#c2:�l��ڬ�6�}C�OX���^�.'��ه\��5:��CbJ9)L*|}}b��h�C���j�N�R,����y�^���e��ʆ�c��k�9�X	 M|g��
nu���y�����A�?l�Q�^��\Y2u������=6��ʑXܑE������vw}3[G���U���\�ZR\�9�j��Ď��_����`v�do�h�NV��:P\\R�Yri��~�V8,�Xh�7H�T/�w���د��(l)a�h�Q�s!:k�-�fe�A��yV��
�B�))����9� s���H&Qթ��3M��g�B��/�R���Xt������!�j�d"��	�N2S|b{<����&{c\j*3���ij8@���	�A��TP��r��$���Ez7w�N��+�6�9+�TP�7`�x���ޅ�U�#uvv6�R��U�^���ڲ�aV���q�������O�L�
����&����Y��;dz�����O�(&��Imgn��Nt�C	q;Ġ���xmt;70�ۖ�D|�)�|�d+�;��c�75mk����[[X	���с<in|!S�k��;{�}�|k��h�aq��\�PrU����Q#BG3��3Mʞ�"2p�J�j��L�%OS�uJ�c����vb�E}8�:����4G��22н�I8i7���R�57GS-V퇅�C5����+�Lcޝ1���jG������海Eb�^���|��(�*�Qu��E?+c���y�u>Ͱ���ߐ�ޒv��sVF��E);�v��*���.���p>H^7l����t/+!zD�G�l}���Q�2>
��a�cz�oKf�-���N޶��׽j���.��z�����a����m�or�\��LyB�VP!��ۿnF%Ir�/�����;���C2%.���\s�ejCq�޳9�j�3����-��B8;`y/�>��6�M�T���������蠹{I�+}����J�CԊd::�KS�,r�WQm��lgY�k�;h(7\�}�ޏ*�3j�M���8�8���$�i���,:j��Y;<j�2K�KB�"?8��xHR.�,�(���yO,�h�+�����g=}*E��\�rA �	���_j/�Ş����QS�j�5b�]���4��/}7��>V�p_s��D���2��4�@}!I|� �Q#ǱUR��_]g��=�E�&.�v��$�=�׷�������.�il|e��y	�b.����u�D�N��9��x�6vϯ�4���rrr�RR��N��c��T༛@>��0?S�>܈'�)���p���V��̜5���:��켏K��
�"mU�Ǒs�avz��f���=��=?�낣W���6$�E�孛ە�K�ҳ&�N��z�\�&�.�:���}��T��)��-�iN����#�|A����k�N+Z��3���ǰ���;.S���G�8��$����q�6<��L�[����p�t2�>��|rQQ�S77�)g����T��c����4K�ٔP�	4��4L�as�+#�@�К���r+����7�D| 5����6]�r�SZ��)�M�l<=u���68��6ihZ���[�:x�O��ZB.a>�Ɍ!x�ū�UF�?�Wχ+Y�z|q'.�u<(z�्MJJ*�v)�n[辤�xȬVX002��ly5�w�u �,j���'ʴ��I���� ��_<��^��&�sY8&�K6�S
����ċ���l��I8m-�$*�n�!�@��-���
L�����"�_�fM������P���.�/��D�AP�E8�);e���!D��5�9�n����7�Qÿ��F��8A��\w��k��Ri��#����Ś��)[�B�T+Q\&Sab+壼��e��ι�n���w�B���v��s�ۿv+}����?Џ@,�WF��}3�b<��ϛlq����6��8��g�$��Qj�h2r��Q�Y�P!�BXճ" j%�XG��8*�� r�̂[���j8����}��W��P�{�P��ޖ2`�A�7��L<�o���I�,��w�aN7a�v�7�˝=g���(Uݶ�����y=ޤ�7h(y�MF�$�Fx�Q7�z0q�Cq$��5�w�&��4<�J������]�b��3�#�]i�ۡ���Ն�G�/`������(��3Ieī���<���^��q��h�\ӭ��/���+����_{}��2��)��}C��E��ݍ��0_Z�a�4��y�\Y�X����L�N�UTT����V�'rx�Ƽ�O��!u�	�<�
B%Ǘ���>�kǒzt�� ʧ��IbX;`NZ �ą��MɅ{����2-�GU��g>��ʒ#�(�]Y}�.����L�%$sPS
�|p�ԐD� �M�e���/���ĂJⳀ;S'�>�9�� �P��}���ǵsm� 'ܕ/�+%��3�+۔41jy�O-�7$e�N����y���%�E�S�g���C�	�����@3tA�}��͍6͞�|����A�~$F���(:T�d�e�L|��M����	m��i�^��?��ݹSGQ�!S��g3�:������X���.hO�o�p�[c1سu����WL\�8Yʢ���b�?�	ND�Ql>�:jX��
q��?���%����#�W)���W^�i�w�P�WZ
�d�5���J|�ŭ�QB�� .~8	���A���6��D�M�Zc�ޔ�Lx�vґ�6S�&�_0F�+1d4�q����,�	u�P��}��� ��5-M�6m�7Lk��1%,b�w�'���3���zF�^��L���&V?��ץ�ｦ����=4��m��N���I�����g�������ܐ��UF8z�-���V�E�Xi�	IU[��M��;;�5F��۞��QĶ���ok}��������.�b{�,9����{�v���,�%�Dh�^��ib����CӸ�3������$ciy�6���P*����O��t�[\��������<(���D��m������h�ֹvy ���<�Se�594�4X���C�Dͤ���,�)HT���Iw���}`5Q�?�=B�U	j|�/f���^��q�A�Sl��p7+�_�4;-id٬)G�
"}�A+<{� ~��as^�������8��ͅo��6ܦ�c��G��BW��7�}�J�_J��8o�+ ��,��r0[.P�t��Γ���v�J��(�S��PoZ��"�F�Ϟ��\-�w5��E���F�C�� �':��A������W+&�i����F�bO7L3���*����i��,����>�޽�s��UZ��I�n��[j�ZS�CU�H�	nR�����(X�/��X�k�f!��j��m}R{~�Ph����2�,ږ�!��PvU�*�OG�*Q1l��s�N+�I�������r�$g\h�sYVq�?�@qb�aA�D��ʝcn�|�f�W[�gV$$!]������V�{�Uqw�����]���w�!�c� ����p}�Zlw��锠\� ,hN��4Zt���V�n�'�W�}�	�U�-j����o�t9�1!3X@�
#a��1ٖ�;]�Š�b,�u��z�/�Ď�fA�?~���˽�O_�9f/"�0!zC�C�����j�X�`��O��ڇ��u�,w�]2���j�a�����<:��Yu�ygNa����),���FcxW���{+����jl^�xk�2��ޚ���@�U�umi5
E�gQ>�K���uH4:̯}�-�>�S�m��r���@E���C�zuj�:q�\܉MLA·�9�j��\�=1)���V�
"��<��«K=������L�g#��10��ph9'�.F(�@u4 Fh��Ghhe?Q6��<�����y8�T�5�`�o�|�/Rd�������hz����{������o�+?�a��RBF� �$�k����j%�w�"?�� J4)w���ͥ������g8��l��k�S
'� ��^���W����}O�'��~X7a.5����������脓(��P�Hdhoω�_.�7!0�D�w�jWB��kB���F�ӱ)�����xyq�Ț��<~�Jo��
��	�8G��<�9��oT���7�����:�YC~SD� �����B����m������Lۘ�_�x�@u���Ńm,�˻���!��s��LV����j�c�o��P�cC��`����W�V���n�y�����@��ނ�8%�Q��l�U��j�E�Ǜ�	á�i7�2k//��p������7Y������^��iȲy��Џ��t��:U���}����H(�n=n¿ ���]S�:�%��0>4�/���7i�Wx�TR��뭾�x��K�"���f#
v��_3<Ű������H�!)s���Y\Z���dڀ�|x��y쐼?zz�b�%e[���0�ipg=�����W|�:)魤��M�vl{&5�֡�G�*ax��&�(p�ٓܨ��6��-��/O����N�e��x ���vJ	��{�5���q���"d�æ�mh����k���}�G�������uE5+�Ϯ@N��ЙF�?�8���SA2�X��ɘ6�|�7�Z��!6���g��j~:~f�޸>׵�j�FΏ_�Gӵ�6�r�@<������b��\׾�������R��" P���8<'.���0yC[<��:n�B�/��O�zc�1f;\E�aq�|DrP���j��*DϏ�s��.#L�~DF�;�+]�����j��פd� �3n�ՅøLos?l5�C��5���hnM  ��-�t�oG�x4פ���=^PR=��H�/S�3z�!��*�޴�����;#-�A����^���Ō����\|��¤����`�P��`0�ө�����~�@��3�I#��<�7'��jAɹ��a�d�]z`��� �+a�و���OC�#���vy��fV,w�e�%(i����&*���rz��:C�h'�12r傿�{@�����XJ�~�Vd�h��4#�j��iW�s`VCN[H�K�{<��\��Q��TfV��]�m^��όc��lF�!�9ل NF�5��ԧU��~/Q��������ʱҴ�.��|Rz���5z1�k�����'Y�7o�"�R=�����|_�4��^�+�!i2\��I�����p.9fW�&ط����DOb>��ǓXq�zzH�&��	4x�d������1e�K@M<�E�p�x2utgw�;Ԕ��/�x�5���Cq�{q��`6%^�(�2̜.[���t�ƴ��էO�+��,ر"�b��U����fy������6E�O�����[�9�8����~��}!)��$�M~���hnc�q�v�L4�����p����q�D����Nh�1Ud`ꯧ[py��6Z�� s���m�J������=�����>����6�ΛՃxOˎ�t�+������ҫ�#��ڠ�Ј��w��x<d�DHn��i��g��o+g��m9b���nm���4�����Q,�iba�\�SV	寰��Jb���0���e�zx�+����"8"�M7�5�����s�W6C˽���%P��Ύ��|�9ʸ�����T/����E��=��`�6Ϭ9�
�8 {`��_dAA��Ke���;F��,Ow˅ee�lӯ���I�{v�fFSK+�ʁx�d`�z��}�LM��~�So}���]�l�\�p��C�gW��?�_m�0�}�y舌~�pZ�@������^�^����T�4C�:[P�e�ih��M���݁f�M�ZZ&��X�k]wdQ;����d��4Ѣ��}�͝�ͷF@N���������J�u�l``g҉�ߥ��Pbv������z�� Ը�Y^��Ϋ+��_=���~|{žv�3N�C+�Fڂ�����Q���Ғ��"̎��-n���9�|x���|��H������3x��n�-��*�����T���i���_��D-��w���{5F�=4�4��ض���kT���������Y�6-fU5��9��ן�=o��d�u�4F�!Л~�kH���O����m>�p��-8+��\dl/ʔ�J�~�o/���CԟZm�s�_<�1��0��yZEM^��:�c? �����K�I!�u��#���LRix)��qI��*x��j�T���O^������ȏ���)��u�~u�i����v�d�f[zQ0���q3��v傄"�d��Y��<.���qR�|A[F^7b�?~�D���{�l.7e����t~�?[=�H�O�)�.��,���r?8��^t�p?��;V�{/�4s!`BѰ�j���V"�U��GbQ���k�%o�Y���B�}%a�O7q��Y38�ٗ�qv	\�v������f0�{���ЋY���<�D�b�>GJ�6�������������S<�F*�"��ݝh_�-�x���x����a�5�h��"��`n�Mr�'�MV�c/���^��@��)�6 {Xx��^I�On=6ru���;lY�l}� \�)y����K����<w���)�s�ۘ�-�������}�A�yۢ/���ꂮT�p��x�9�L��@wJ ��d��}�)#n��4�ڃS��=�:�X����r���k����ύ뎁aa�BKo`�~������7d���:eDj=ss�L۲S��BQ��-n�ku㒙��^�s�]�c&�E^W!)S퀽�y�s�5&�'�""w�Ko0��*�$ܑ?���lʴ���mtd���j�Kf��p1���Z}_i�M\Je�w]XX�=�7�J�R��)2I7r��&�;k���H���h�x�'��i~D�[Z�j!����B��F�[� �D�w��e	�'��(�e�jO��6*��+���N��8 Q�&�a��&Ҧ��{ۣ�;��p�u������ԷX�����v������G(�n\�݇��C���k�ϓ��=J�.J�Z��2���d�.bS�b�'����춱��3���k{�v��}ԶY$�$EJc�K7/����N��I�Gu�?���#���R�%
edj�u���㪓��>��ڥmo`���[�ι�B�o����Fq\���T�z�p�t ���Ti�&�7o�u��䄅�9�\[��]���e�ˇ��o��q��nH2�ݎ��܅��f�b��I��C$:�6=!)z�9�s�d��?�܆�W�ܤh%�|����R�Ϳ�.%�R[ØU�����yf�0j������e��j�a�"؋{��}��,膂�` y3���n}m��<����{T�@K�ׯ�5�tb��r��yJ@B^f(1/���B?�Z
�w�V_{r$a׵״ԕ�i�|������a>���Vg�OKN.��G���=%���.>>���J~���ᡴ�Lkk�x0�_AU83�l�O���f���Y]�PXQ��^w~�|@#>^N��#l�����s����3���\L�T+�Hw��z���?���?
�!*���.V����z~d�Sc��9��oOM!�ܬL����vK�P�~Ů�4ZW2�H��jE[ß#虀��ݷ_�T��^H{�l`����k.��_-��"�����|�|y�����<1e�jz`Of�ɮ��,�ͻ	����zv0pߒ6E?��?�P�*���~����~xk����h0�0h ]�s�}��s��ޒ#W�cJ�I���#X��g���R���X�����2Q�
?3�;��pw�#}4&�&3>����sa33���}�"��������Ea2���Uo����l|�Ƃ.��jĊ�@�vG*Ed�os�9�څ�l����d�^p ���g��B���m%o���LZ"�R��u�W~!9�����=����v�Ff�1�So�i7��+�0��6��k����d�W�_*A�i0��O��Nv4羿'm�Ub-\D�Ծ����K�mZy��/ ,�_Td��bj�fxb ��B���^1���Q�h���-XL�%7�)�1��i�������8�l���OOh�\{ ��Sw���ysǀ����Q����gZ^�{��xMT<�<	�-6��'I�;X<��~��\�TY�Mg��Yͨ�J�%�l� �p���$�����)�o������]��D��eK(l���)�&���I���o�L�z}}���	1	��'*�;v��Cܾ��P&�,�9���8�8?}��+U��MF����H��3/�~��f|�&�X�lB@f{�;���;�G�A X��~A����m�).�Źs1:�_c����������ak�ɽ���[�r�\�H�O�}�8�k����ST�a�t�G/]���ĕX�~V�&@g&e��C,�Ȉ�{�Ģ+-Z�|��:W�SW�A?Y�w�J%u����r�G;>��{I�s&8j���jK��&q����ή@��6v�f6f���i|u�mykF�,<(ê�]�4��?�o� ��G�}���gW�Y�I����d.N��:7��:낈�%��`���Q��e%���Tt	.m�z0�Ƃ��ʸ��]旴��G�BJ�I^�����<�޲��mص2-	@?�+��� ���|�{2�|u�>)&
M�`���g�:L}k����-�#�f����k�O�r<�H-��7�Ğ� lU)������TQ
8%�z�x��t�gR���{��}r�4�+KĔ��k�7�$Q�/>�Қ��9W�告����~�UC�	{$��L�%=��ߙ��.��M��Գ���Q����U�@ݙ;:����a���T���B=���n�����.K���[{��nb��Ζ8�� /5�7�8g'��_Zc�L��.#X.6$��XV�Gɽ����?['U�
n:̫.1���q�(q�ynz���Tc�����!���R�ѯ4��	w��:�P�L�:w�(<�U��\!��/�R���P K�G���!an��C�XCJv�I���k���E~e9���B/uǸ��yM?��L�	pq�\Z�aJs�u-C��j�N�1�C��b�M�6K.�Ő�O���Zc�5l�)�T�œ;]��P�D{�y�y5�2w�W�Az��گ��pF/ʜ�X����@����E��u2X~�}ł���h7����IfM��7��<�/G��6$�
E����<y�~��%�׹g�<��/&���#���X�i�!Z�BJ �Ęť��߰�r)�-�뿅t>`Gↁֻ���1^ab�����K�	���|l,���7tŸb�k3؋�F����س4��G���=<�'�OK��ūR��Ox��rP���ǝr�g�{��;<m�k�����ȶg߾"jG29/Қ�I7a�r1b�ݜ����ZN�Ҫ��ޓ��\vm����),��nR�/q@qd��4H�	�f'�z�'F\���TX�q�2oy�����JZA!�
����ի�H���W����/��r�'J+���C��RcH(�u�K[<e!ca��e۞����ãǱFsΗ�-�Ce����q��+��p����5��u��u�8�w��l�����o:d�_�<��y����4�W5p%*3�\�7聍�w/�|�g�άύ��xq}}�����N@'Ͱ- �8zaƓ?�����~Hn,5���!XcY��aW˸H��-���b:15,wŭsE�}|?�),'�*v�w��	K�����Ǖ�l���T$��dq�2�~�VV��ONK_''��uz�X_�*:����a�m!?#�z�q3���5���G��q��k��6�Ć���I1��O��$��G�`Ii�?3P�����_mX��&���F�?�bG{����"u��N��@r��q�!h��������f�r��G,< �=�g��ma�3�a�B�;�J$�z�^������\��=Kr/x���>a ����xo�}��*^��٭'���ڔ(��G2���"����&0}�a�i���x�4�[�3�f���_�7w+�P�>x[S=y�
�7�گ<�!˃�i�n����F��$\0%�&%2����ª܂ZG���g�$��p%��cVI5{ ��+g�1m���#
�O3pYUFXW�Ͼ�=�X��4���{�чxZ�ƒ�hƭzh�I�es�&�l����ݠW���^�N�2J��)Lw�+��K��r������_�]�W�`�;O���-�3U��~4��X��b�M�f���bm��BR�<�[9g�L��r�/˂������MQ���r4�ť����J�}k���o/����õ�vi��?	�� �2C<t��a�j&��~Á��-�d�kݗ!E�<􄆪��d9m������+*�:��V>�����Y�Щ�Tϑ��9hd�7@q-��7Y/��_-�Xr�Z��]:,GFb��b��oS�\r�Vf��v��p�x(��c�r����JC�o��/9Efݻ�������yy��#���7������^o��L�w'�O��"�T���*�G����
�C�'��F��B�b,j�|:�#N]3#�ĵ����=��ψmӯ6��\��X�kt�I�9�~���(5�N7a?{9DuЗ�lX�TY0&��	~��Ux��ֽ7&�0C6�UY��Wܼ��6O[#dd�����	�rZ(_7k�ÝD�;n;���K)��B ��6�[=Eg�h��	��3Ew�o�o�Q$�d�#��v��g���/�����B��̀��z"���d*����5��r�O���Ar��>�h��n�����+znY��[LJ䕺x�*�/��HW�!M+;C��w��y"��@vl9�+�Z�]t���,��:�i�t�T��%hT�ц����<޻t�T0Y
�H�-��\�8�$I/��j�l1K�����'�.�8�8D1>���޳��~>�`hb��;�'�៉w*���Q�30:�#�P���
��p5�Θ�/]0��p�:C`M�����2���v	��ω}����)U��nR�Q�&����T}2Q�ր�X�%�� A����k:O9F�[�d��$�-�u������7x�a�O���l��t���	����E��'��}p>�+�SA�-Q	���:�Q��{���gn[�OD9e�4�@N�-��7����l�r&���݃��q�_�����Nm5���)QzR�z���q��v����%��Ǖkq�Ŗ���u�����Y�Ý���mW;8|�Uk�r?`J/����t�5�!��9�A��=R���jϾ�8�c�ӗ�;s~p:��V�M+;[�����Q�4�5�>�͑�d�ؘ�����BLOW�a�z����r�eѣ�a�����;�B���/�_Ƴ8���|��K�`�a�p+��C5�D�n,9ԋV�����6"E7� �� �|W�e8c��\�F��-�Q��T��&,4ڗ���F�n2׶�w���Dqd��cߺܟ��u�L��90S�w0_׮���e`ް?c>_�2��$��FL�ۺ���I4����a�/���{}UB���$�.\�B�B�vm.4b�nUd7�A�w����In^���p�c�4/#&����LLM�s�*��+m�0VQݡ�b�l�{�y#p�����U&kN���Z.[��+h�&��P�KK �Bհ|��[`�r_�[^>� ��13[\�G�����3�5�qB��������^�x�|���0��z�98�X:�RE�,0b0t�����+;<^ݞ������Q�%mW�A���=�a�+��&ey�T�pL��uj�m�t�]����`F �������ʠ-�_-AE����I���!��ꝫG��k���َ�%p5��9��6��'
��{8��{u�����)�^�TNӰ��Y�݋��:	1�ޚ*9~\��8�8)Ҹԓx*��ah&T20xv��o��l.�ײr�����`od8�����ug~75a5a�~��^5[�#h���Vk�C�p������8M����ұ���`c����z-"��-�)+b��Q��H�	py��A�ok�:6_B�8],>�l�<W���Z�5}��7n�u�(��**�Y�S
�̚��sܗ�G^B�}CVL��&@f:I�Š�#�� �w����Q_��P-�-�D�v>��Bι�h�vx��FZ´v��J���w��9����!q�N1����d�ɖm�6��{l���}������/����^n�Q}�4�����+�M���ye%^|8I��	[��.J˳C5����fdD|Ik���dTdJ�J�E��~c�g�$�rHZ|I=O�@%���ճ��`����d�u={���Õ���k:K���w<7G]��FK�Xx�L�b#w^iLJMH���G,�x�(�/��3���jLC`�Tv�ElAS=K,XA%me�۩w[�ɇ󉊮�/�Y�ŦG��%�yg��@�������vP��ᡗ"�i��Ɩ�f�Y�! �u�Yd;ē� �;�]py��~UN�]�F�n���MM"H$�@�C��|��L��
'�}4��V�������ʯmeQ�7,x$���kYٝ_�J�%,�(yI���|�Da��;�x�G���Y;�$~"�. \��7�#�=��J�'�]㧷���G�ͦ�q7��R�O�n��|j���C�ƣE�dq�\���'�������O.�rum�I���첞��T���"�Ăr��H�$rթ��Y�!����I��V$2
���G��T�YOʸE��w`��h�=X�-��հ��Ų7����ql��0�T(s��q%#���>����[\�M{����>��Q�6��<Ii	p��7&
��[nh\c
[nk�����^!�~��s��J�MN���� �!�&����R���u���	��T�_8=�:^�\����i�a�S�=�MG�N�����ݫ�w����Y�M��<�vO�x���}=�������!�*6*
��g'ڰ�����$�ʶ�sz�}���_��	���(�J�._�ז��~+vCn�z��_�D��Bj�2|+rA]�ƃ�Z�r�N@�>OaG��H����`F�'D�cV��zv\6T��E���t�ms~F�t�=DI9x�ۘ�Y;��1�l�vh���l���D�:�#su�D���,������Z�*�	���X�e�T��l����'����ԑnCp��U�~��WF�_��6ˌ->&�M��/[�,pi*--�U���Ը	L��\lm0=��t(�Դ>L�b�Ӹ��&){�O����6u�>X�SXޔ��������?�S8�tf�S<e��������@�3�ג?)�ѝ��o6	=y����x�'�����ϧk|���'���C"��##;��qSMyyy��1W��6�e�Sl�6�1|׬c.*���:����-�D,�t��> .�����S���'��5̜]���d��x���c�u5���+��Ë��EI��~n&k�X�k/~��Q9�6�3�F���M��T{���ԤGC�]�^Z�r�;~�Rܣ�ǐ���_7�aċ�X�j��S7na�Mvwy�w|�s�>�[�����Ebff�����őL�&)�շ5� ��f�<h	��,&`��Y9��=���x~y��-�y��^F�y!J�:���>(7<r*���H��������d0% ��,�pC���P�F/�f��+��a��z_��&pP��U�qY�I�/��������J����c4�93a~�}�Ō;8���;�p�/z�M�&�uч^�������>����{AsːG)�y��۷m��x*�**.{bZ::�#0����q�rL�] _^�_�6�_��ډ���T����ߊ��qb&��g��W��F2��k�#R�h����?��8�E��y�i^�L6�BlA�y�<�}�K�[�Z�ƨ2�'�pE�Y�^탆�	��y��J�?m��ף�OXG��^�F�6C��ֳzEEA!a ��>�J����9��i��PkO�AрU�UT���(#.#�Zw˙��%G4R��y#G01�"n�b�?h3�Jɰ�v;�ִ��=֍�.3�G������i=�x݋v�=>��ݶRv&�2`��g�}⫧]����F�8�J�u;J��$�.��2=-2)�g9V֩u�3����GI����L�o�\�8�u�I��.����\��m��M���g~w��d�E%d��dڀ)�M%����t> �S�l�������@,#
NdŸ���v<�d*�qQ��M#���-k��Wd\��O&�/���<.Z"RW�����F��� �W][��Wx���e$H'�T
�s����#�v%c�pct���=|��`�����Wƃ}'�y>t����,���n��b�o�ESc�d�|�M�z&�oii�Kw�=a%9�Û"~{(����K���(ْ��]{a�G^�ˌ��ͅGhC-��@��ˌ}Ï�`^��^���H�N�O�>���9�l�qC!��~'����"��;:Q�zW�r�ܼ�#�����E����K#b�`D�'Q�����Vx��Шk�Q�N�������H�;�r��4|�a�#pB�xE+�����o�*�<���_���⋷^�������XT�/�;{���R0��D����\�k�T�E,����s���:�L��YƯv���m�8������ѧ(���$+% ��;�CڹSr?��mo�G􄰲�6?�߭Ơʾea�'|���>��[�q#o�+���no�)R��O�~,� 7�A}���ea������o9���3����MO�����bPt��B����}�3�؉Ա��5ރ�9�$���u�CZ֒���e��q�t�=z���}�UQ��/�8j��G�|^�C������7�^d����I��JN7_P! RT���$����$�L��Ҹo��\)K�������6R�y9yK���֗��4�Y�3Q	ɹy�kV�T�eX�[�?L#!��(��t#��ݍt��t#  -�1RCH���R��!�0�������</x�u1{�����Z�0z����D�	0g��S��xTN/��sO���_���%��_mcJԑ���X�N�a��ٲ��HhX2��I��@�) �)}[�AFۭ��kvf.!���Cf��ٮ\��t���ɗޚ gL��&u��Z�q��,\�����mi�B�>��Ij�H-�(�<�rF�Z��aj[�Tڗ�D�S��;�F<F��I���Gp6a�A)NO~oV�����Z�t��Ѳ��>�vP���;!��)}���Ǡ�A��D�cǏ�;��0���%����WrC�����$��X�xM#P���ޑ��m��0�+Y��g�`M�}���-6���H�B��}A���.�)�.�1µ���$�>Z����%e���%���BA�丂^�T����
"�yo��YܢN�<���rÔ&�O��s��{�fS�}F8� �$-&ZD(���M��蝄j+%�w��N�#���I�l���0>���Z��=�(�_s��~ �d��2�C#��sh��?�T+b��_q���Bl�r�I))6�}7�K&��=AZ:	S|�!�6�" ؝lO����V���Nm*�F��P"�����D�xla�naI���Z_2��D��CJf�}�6�/M2={��h+���P��wgdA�jY��{tV������S�\_�ם$�[_Κ�]LⲆ�����ҫ{����Aǫ���Vm�R�{�%
�n��w�w4�������b��wM�L�h�8�g��"M�8�ӠT�	�*�v߹�UZ�<Cn�uy��wa��B�{���Il��т�q���6��Zoy~)������/:ӊ ��w��X���dX(�}�w>?
�Γ xq�����uH*�P$6�B��tR׹�v�*S_�����I�D�>�����R���3��r%�6Ɲ�@�KS���"������ə���-�k�P#<<>p���ycEVX�#>��pk2ʤ��L~�Qo4^�v��� �����ʬbt���²�`)��N�Cx�kvO�lcy��@�k0	�C��Vt�H=v\���CK=�0v�jJ0���k��+��	ӂ��2ؘ�~�D!�n4#��6��;&!\vĈd�!gp��#V(�h�5��0���Hz��'B3�+r�F_��>9������� ��-Δ�W�����ǅ	��N���������	�p�f[��&�T�;�_~�x��;���3j'�������Lac�U�ͼ�}N �+mϏu͖��A����Rm3�B܄*�Ǎe¹�e�o717?�>�_����c����C
@V�K��|D#S�̌��J���3��`��._�W폞-����nX��D���'���\�n��bͻ�?��5�?�[.*h�t��֖-odK�)�%-�:lJ�6��Ĵ���4�g�薪L�I<��}�B�A��s^�Zk�zE�C���0��/~�p�z�V�*��n�S��¬�J�Q�����Ќ��!�p����ö���5�4�%5~F�.ܧ��ݏ���ܰ/�+����ݜuRSU3hi��B�v���ym!~��Cu�X6���'n����6iPϽg,|�E+�WZy9C��f�<��x�0nQģ[;__��Kf�������&��Ć88��&��`�D�6����5�ܰ���Ү�������h�p+������1`��[ʡ��MwY�SK8�G�xKZ��J���	Ji��oC��Xp܀ ���#�2^�t��V��[3Z|m��NҠ�d�(T �z�;���;d����h����שWֵ	0:U�5��o�����KzLo[N/�5F�`棵����E���Gy��y���E�'&����0/�U�_�	���޿�:T���,a�L┽:-Ҷ�HIK#u�hE��8>Ͻ�@_� ��GT}P@ �2{**��b��'����/����&#�a��6�ؓ�:��tP�ն���U_�x�6N?f%���hXz�bL�\ŷk��bǁ���T�˷��f��������ߛ5�����pt�$�_J;l'_��%E⓾l|w�x�&z}+�;4�s�\ƿ��=ƛ_myR��P����T��?ko9�~
�ǎ�b{S���FE�Ђ�f�JKK�W���`���}]g(��'����A&�{��י�i؀��d����:�1��:V�2��S�Db�d�	��v�[(yg��J
�t-���'���wD���Z2��|":��>�����Qg��6*d[�'�Hg��PS��O�^Ćap��� Y��b�^K�䷟d�Eք������VA��e��G}��O%%��4y����?$�g5��Veى����gi���t>Q�cTQU;�Hb�� ��-'㐤���|*$B�/��<��e���d$RL!E�I=���pe6�wR@ޑ��a�p���[��
}�$��o����5k��@���_��Q�p���0{�*�Q"aH-{-�T�K�=K�#�����%z^uj}��u�����ЖE,���3dqc/)�^�Q�7�;��߉���������.���N:��^�f�G BO;X����]��./�v�h��soP����'�;��lo�d��:��$	qh�y��L�	����?H�o�ۑ6��x��Rc��ǃ���G>=gq	-��{��A����ނ�[jē� �T�ӣ6�����q�J�FX��ף��fU:���?��w�sr$��]��d�B���J9R�?�x�k����`+�������ǌW��`�j�Q��a�Ɣ�Y���[��8J�O�� ކ]��ԢR���7E����~2+�������I�Nr��O~u���O��ێS��IQ�[�E!fs��<�㎊���H3){��&�����L���x��܉��>�	$}�����O�1D�ͨ�IU���zW��{�����2u��]O3��u.I.Þ��+�KPH^͸�q������8�Je�9e�d�����j�[��Z]�ͯzS^��g�F-:���U�X�a����Sfp����
=AYٔ	7COp��W�d,JJ���r�T��8����:�WFc\���sr��oz�MY;?��L���{��u�7��+��L�3�C��G�<����寒򵎣�� ���w�Y������w{�)�GK���R�D� 8_`�c��Q�o[��r)8��M@�3�������»���� t� 7���1�������fB���Q�����@x�0�߳��|.�,hL�`���ME�B�	P��{w���V�j�t�X�j�c6�[�?|��֍\�H9�Vs=�	�	���BM/���큖�;h?`81VaTZW��M����T��.�ݒD(��0�盰�N���X�>R�Ѱ��-�6U3�b�@�*R=e�<���~]���05��wFvw\k��2�5k��V�L$��~@7����j�]�y������Y��������"�66X�&���MV+�u�L�2��k�Q��"�6vv�����@(�e?Q	��񉐭��J���fS2$�eÝU����p�����q��k0���	ц]�����<1E��{n�	��Z��AP�s{� �L=�b���rW�<��~����>/�u�3о;9���3.�:^�d�$��+�9��!*��4�Iԫa#�k<����7��j0��R�:C����7�}�X�FF�$���f���.a0?�Z�W��
Y&��3/���jQ�KR��'�Mq�~1�}Y�`'�OX��Py`������2��/EC���W#������@VG�5y{�j��[<��}4yQ,+�_��L�;˦*���{(7e�hODc�R	���P"�O�!�|+`�7h��o�w�!=���.s�4vǄ�!ò��(��OL��2Ѯ{.a���R}���fy;2ݴ��e��[��l_��b ������D)/�e6�e��zT���آe%���q@Q���I�f�WQ��?ߵǔ���r���$%���9�k��V�d�w !߻�)@�����~���U����m���o���fgz��7��3��Z���"qta�RR��I###t�H����~U����'!)����������{�)>&�᝹:c�FN|2y�3p�z06	����"����B1̒y|��*�H�}���o�X�d���6��Ï˥��Wo�zuT{we���<����d��gJ:Q��'�/�"^�kf�N�v�c�+~���|*����^<l����v���.���m����dz1��Oѳ�'���]V�,�\���U��J��$�W3��5��3E��dOP���x�sV)�Ϥ$0;�yn�(C!�Yp�WN�t��=
*8|u�<픤o� �y�:��Ȩwa_�!^,�׉kp� ������ry�8��%�5�
���\:t�����R)Ļ�~�&�bT�L�V�"��_^h]d袞�Iv�S��B��Z_�2��#�>א01�mX�k���g�=+�<�p,��E;��@��w�����¸�/����I�O����k:�H�!�xZɀ��|�@�\SQ �lmm%db-�������|��\X ���f[�Fyr������#��V?�Lv�@o��������݆��a�{JL�tFz� ��Lg[�'����NN���M/��k��2�b�7t�h����,�E��S6��Z]����<klP�>v{�8`��=��O�E}rp�n�_�S��{�j����J�/B�iUu5؇��p$@�m-���I�)+v�=�X��Z�'�0O2s8���D�K���ۓ�m$�*�����F��O_z�O��\�Q��DI �* "�4H ��qɳy?^���]!C����py�uǽ���%߰^!QɄ��[[�)��ɓ�I�����Z����~5��4G�j3,��t�t�Y��O�F+������㟭k��cSS����a�p[q?��D3����+��Zfe�+�Z�fD�w6�s�`�a�[z<#�:�����
o��G�_�����G��#�Q�a�m�b'����%#�F�1�]*�)����A��'�!����0�����`۹)�����������7�!����]���*\h�U�)A�ɻ/e����l/�׫�����@<?#EUE�9�jaar�yy2�� --X�P�Z__���.�.��Kk����{�臾��x(|A��6�B���e��{���Ĥ���-!���G&��m/�_E���u��;�c`q�LM=�j��	�L����� K�/�n����S�s�ڔ����O��7�*$�j�!d��	�w���aL��'��,����C���O��c	5eN�R��D+��-�3%u��WM�\�8�F:�)z�zwjy1<����U)�U��9�o�����~a�{���y#��y�=�~�'����s��w��d�2V�9Lw���^Q $L-T����]���L�j�vޭ9)��^�P�Y;R^=
���:l���z������I��ex^75���~�Jb���������<0�E��O��{��꥚���ib\������;*�g,��\���ed +X����.�5�r�W������G�6��������/�R�G��~ɮ_�sx����0���d��r�@�6g���0b�h9����c`*�],��0�����3t]��#{w�'Gb����;��-k[eb#�4����\�A���gE�x��%�j��N\�������RM!f��&@��7�<�$pK��b��-�@xM�`V�0���r���崸�R�SO�1���y+o{��)K�����O�%�Nm�+E�3\dW�kΖ�i�=���=�n
��9d��R�i�jJ�r��Na�4��U���"4�#DN��9�#�krr=Fee�#�9NAA�Q��`Gb��L��ш4;<$d��#@�	���b	�}�����e���1�g2�)T�L��HRRk;'��r�Zh�0��<<2���9﫩����㽰;\ � pѦzu7��{m8����w�I0��_Ow6�=ǎ�/�l��F��F2M��p��^�ojf�^����mc�� 	���ڈ��F ��Xr����!��Px�/^�m�;�r�ca ^�� �<a�,���f�m��+ٴ��b�yMW>�xM{��N��HĐ$Y�O+��ɜ5��T���	�.~��S<t�%퍤���}����6_xmooW��3�AX�Ɔ��V�i>[y����v��7<|<Ai����7�4�h���Oϲp��jK��@��u���!;+�/f�/9������=��oE���>��ND!66�c�`pYX�-����.©�T��[@G\�d��S:F���}]����U�%2�5��W�:�`+�w/[ـ_�
'��G2�I�����͕�V�F�%b�Svo�agD$!a�0l����ޗ�L�z�$
��<\�{���!mԩ�F�93��|����T8�V{��C�]/��?۰�T���Q��B�LYYa��+�B�jy����T����M�G�	�#��֝��Zm��p�9�#�>G�wn��a,r�bs�X!#�=>�)�m@��c����%��B�����a� ���>�����)7��3���n�潕�k<�6���]+ߦ��O�Z��55�8�)Ē�l2��P��m7mG7��Z�Q�ЅfGRIIɲ��ψ�'E\D;�,b7��F���u��5fTy�^ASJ[
���]cϢą����5�9 �׭[�ݲE�g�)>dgZO��V�s=s~��_L�T�����w�K��R1=^DMB�1` ա��:SZ���S%%�|ji�z'�ak�U��}}F��el��;�"�D�/SI�~�-�������,���KD�j�}���
�ʕ��5�x���qy�O&�	k �v���g#��ԯvK�0O߻g���x��(Tl�U.O��W��c<{�����ASzG;Q�8�Jdo�}}�=���3��W����>��� T7���f�&`Q�/�]��"���8T�* {�E���Gc�f�z�CO/�>xv��/��8�{�ZUt�Ҍ&{:4:�ibb�>�TY����|Y���6*���-O�p�wm+;;��EC.�����45[UU�< ��yx��%��Dd�\��" l��E˙oqs3��R�M�K�E��pB��qo����s<tr6gz*���=�{����Nm.��W�L
#�Ap�D�1��&�H������㚏�1�gQ�p���Y���W����ܾ�Tl<C5�}�
�ׯ�(ʍ��C}�GU�|v���ztG�]f���i\O0�"���6�`�KLW�Qn�βC�綌sn��M!O,\�JDWk��R�S&��-�7��>hu�=�[�Y��&�ޯt�ȷ��ҺNgf���X1�s[J=[j5/̆� a�0���� ;�Y<X��8��ώ����T��B�;+T�[�`�-â�&6Z�"gqf�>������a�������Y�p��� R"ù+5c����c8�&A.�C8��Y�_��+�<�M�!�����@�p?�d)��.��v���������"N����j"�]�⌊���;;���I��|��ݩ������h���SWG����5`��Ğ:/|���	�;�k��#�3�(_@��B�@�u�����Lx��nq,y?��ο=(��6��iJ4�0�dp�.��Gk��\Ȇ����,ߣ���ӗ�o�L�n�Ok_�/[��4$ y�0�NǃZ�xR�������ӊ�f�.'!�{V������Kl������W�+�3��T�;/�魥X(�s7�yl����������ؖ�ص���,���n�w~2��U�����cXHt���
���Bd]uף� ���p�h�D�_B�V��m3[����OԎ�Q��������X��{�7�r�����i$����=Q������D�Ǜ�+D�f���;�lV�L�
m�D:xV'2�V�W���WC�����{�w���eb�/�������,y�0O��1h�Dʟy�(o��C��M���S����p�0��nQU�!pR�3f�8$?S �Y���_+�nIlf�o��B�"|5c(���_'o�aJ嶚8�N�9ԏ:@>2���(�鷰�8�z�����[m�7}�cr%=��k����Ӣk|II)F]�!d,���w�+�at�M�s�.2��5���VN` <t�pi��soមk[0����߫���ҧ�_�/1Z�����K
�X�����!�@~zs;Y�]Jŝ�#G��������i��C ��TTT����WR�'
���D����k+|&��L��f���M�ϵ�8�ͯ�04�Z�����l�m�x�M�l�/��^fe������;�e�\ާ�;}���z���i��zB���?�O��z O��Wi!�i�}V�c�8V]九-�1�_'i�Lj}CA��!�;� �}]%ů�\�Y�=3��9��n�j����Q]�*�����G�}�F9C��q }���T.AF�'ȃyڃ�p�_�F'���O׮���Y�r-�vҠ|�3z��&,%������J[3�IVN�8��b�ޱHh}��n��dG�u�7�+}h'`&��հ���SA��c�R#������Z�@\�&�g��F�c�[;lv�Uƾ�_ 4(�B�oY&����F�:��ޖ6�ܖ7E�܇:�M=9�ȏ���`�GL���T�9tI)��M.����w&���F���nM�u����x���gAPWbA�e�3_�d[�t\��O�c0�y��ɬ��T���g�j�M���Z�P�������Y������X�`kW����Ŵ=��v�^�9�z���u�l�R�^ژ�����%�U҈��d�#�q���n,��oP��G��ƍ�����j���Eg�n�<aŕ� y����c� `���v,���2����&���{.K�E��q��'F���2��8L> �p'*8LqN���1�*5g_Î���<��}[���
����,��=x��1P�&eb���[y������`{H���ac#L7����'��饈>����.�XTi���Sצg96yz�ƓP���[Խ�>o֯{�`pi_�#
��j�����\ScRXt��6�s�=���$۾�f�8j��SƸľe3�F��Η�S�Ь���"q%�?�@yE��b�B5 4O���IBϥ�Y��刯`����{���U���� �F���t���/l�J�قf�^��s��2�L]��H����/o�t��|-���(L������дq�^��4�U�?J�gy*�μ�}`�W�|5zKmcbc�Ng�ĩ��) {���p�r�i^��:�=��9� ��IJ�ZQ=lԩ�<��>�pʯ1'�b���x1TSF�O�3��)��}�kОM�����R�?��'/t�r��7Ęo���S\�ש ��E{�ԯ~
{�����w�@���G�2��N8X�:X�"���'6vKO~���U�۝�d�^�����)�.�d4�o��/��ܖ��'�^0bE��e�[��fl�!H���7�ӏ�[���z:n5��7M��H�r�vk��;�����{��� 'Veoo�����a�_O%&|�9- ({�;��^�v<*��{�Z�
S=����ݓ)���n,������Y�ۻO|"���AE�WB!ɇ�h��#��w���c�ںl_Ӻ�m�R׶��@?�ig��%G�X��U�pG����ZK���#+?~Q��S.� ���AS q9.dH�����H���ݛ�o���|���@p�,I�{)O�?DN���8�I�ox_8�0�=w7G�eevoM���wM�x7>�W�<�=�Y�������b��'�grl�,2(�3��::����c"��:<�yF�C���o�0]�!ߟ�\��	=���!6G�/�rFq��Oh�Z���a��TG��g9sT���[��9��Ɍ��*�rm�tC&��z�[���a`����	�q�Q�P��)���|�k��{�p�6�tg�z�����+�`>pw}�
�z��gNO�z-A����>��HtTvR-�n�� �j���Ĥ���:���m�ٖH�~��8(���'Se
R��Fz�e(-ZR[$�YP��`T�I%�u3P>Uu�2,��xb�_P$��\���U�A�N}����&�/�>�a�Y	:*��Yy����kۛG���(�¼������۷��JY]�l�9��h�|f��&��Y6�2�wq�8���ĚK�"\&���ߩ�^�������=*�u��N�E]�E�@�����ͽ%>'�FVo|�U�{��o/m<ݲ�_�Ϩl@|�2#��yĊ�v�N��!���:���O�Nt�4���Z�\����wkFB�Н���=�;�t�C���E�C�����������:mtz�Ɖ{���mh'���C�\7��Aq��wؐ�������;5���y�\D�?G�kQ!�޻Ab�6���j, t4U5	�(h���_���	�pHߺ�1����	��Խj�b8r����+z2�GEA�p�H����s�Xs]��}�gR�mPG��m��s�n�B�������ϟ�m���9�op��$.�y����ָ坠L4�Fx�e9X�F�hq�ӈ��vɴL7%�v�/Ci�� �~>�-:t�^d�Q�HS��[ʑݧ������_��B�8��i����Ȍp�黿��^`���N�4�VR��U�#ď���8<�)+�vIe�O}=�q��8,���A��#�#��V`וM�xH+#����A�R��z����y��L�Ċ��]4x�9��ږ���uG�E�ތVg�7��8���$ r�螯?{'��6�|;[�cP.��(��h��/�j�oku��
d�T�}����m�����3���I/M�{Tz��)�?� ��3�Q�-�Ɵ�A2���i�
� z��)����PMOg��&I�a[/��_��g�|[,������p�.6!�Ch���x ���D�`����B��cߧ��'s!O�{[kʩ�:ɞ�=/	\���vJ�����M��}b����z���ug@?�NB�ރi!�ߖ�U���<g���v:���/�m�݌I&�u��充[|��0)�4��(�~LП%Ŏ5��F&?DxG
Lo������].{p���V���WٟxcX�j�ƝTQ��b� �П�X3%�V �3�8�&<Zk�D�,���l�uT�{rd�DY�� {V������2���|N]�k8�u�(*��[#�����zqj�&��a2�y����isr��W���Ϗ)P�1e�U�����g/w�?����LR��(���2d�����C��_2�Q��T0J	w�h¼������~�x�v=24�r��EC{�����w.��{�P��������+�$���Y���ӎgY�:>��ue��¶1՛1�"�^���%\~Ad"�7]#�ȭ(���	1��~ݴ;�
�ZI����5��]E� ��]'6_X�AY�=�|U0��d��:���݀��i5O2��O���[NE�ZY*8׎��/�:��a�
����WЀ������[�z�O�SLI�w�}B����c44vx닐r2/�Z	5�*�^R)~����~�����R�=�G)q���o����{���=*$��_5i"�7�-%goܗ����lr�KN�����Z ȗ����t6M&���) Dǰ�U8ER�-�`�ߠ��񫷟o�m�g�Q�2ӳ���8C@�AA�@
z��H(s�Q�W0Ц��	He�� ű��BU$�Z֚��U@���_<���p{�(���N�ޅ�CKwO3�G*�1W5���A�&E�������)�������kL>�D�,5&��z�{�-6�^�>YC2�w���,�×[eP�mfoǢ�
1Bd��:��?���~L�OKVnؤ�U�E]���܃m+s�0��L�<�����3&�7�i������Ͼ�x^����j�&k]���|��>$h�+y~мS�qp*����T�@�m0:JЇ��2���[��)�kM~���B���yG�M���M#�����B���(٭-�ɋb�e-U?�{%���V��\�.=;��m�����2~�T��~<��L$�g\8���Z^�69L�M��c�B�I�]#��!m#�σ��)3_����vE�lk����q8س��jV{�\ʱ2��+��x�.��������K{�Iar�ĝA��B��1���l�_H�+�ф�곲^=1b�`�c��_������6� ��/X>�V��Uv��-o�x"4����4���&)3n��(d��B�z5�>s�za-�n���&gq?<�yI ���ɳ�#W�H}v��p�V��i�W�_}���99��n������tϭ�I�{�~��t%+{P�u�V/M�t��4��w�������S�ᢹ��b�4,�S��^����n7�鵫�R!��?��M�|���Jm�Rf06���{C�s�4iD��=d�6�|�sص�T|f�Yh�ޒf��K�+ف��|�{�O5ܡ"�?uv.�߼>h7��p�Jr8�Q���<��$����i�7���_��J�E�ռ��c<�	Y��V�H?6��5� 4|�$s��X� U��#W
�)c_t��8I"vū� ��G�XM�쇮Qoh��\k	���;��Q�.���@��.d�2�߯l3���e�����UkM3*F˸����`��wΥ]@����G��;����o�Lw�������v�k�I!�1���;ˊ\�hS��j��<,�R�p�N�e��Ƈ��˖R�0��!��}��Q$��[���Z�y��ҭ�8�r}����0��mʤ�@y�Q�/Q� ���q��c;�)�9>b�gP����މq��
C�l~��d���d�i�6��W�=����m��c���Ο>|f��ܬ����_���7��kDav�)ᵅ���g��BBdzN���h�ke#�7����m�\c����F)��g��WU�(�'��:��+;@4��QK>�[^�d�Ur'�l,�N���mp9iߗ�c!�^lc���E:��D0u��@<eS!j�o�0L� h̀c��_91���	w\��  ��Y�H��z='�ZH��n��|Oh�`nr�yr��^�nHҐ����W��*^A`O�l�Ƕ,�pCyEMQ ���~��5�կ~�Q\��[� <!^��a�y��|y��)�b.�.-��"?���%�e���z��� 5���V;{~*8���
FBW[��S=@�3J'���U�	��}��YZ����0w��l$t�y�q�b�>�B�@��X��+�m��}]T��M)X��K���r���h��|���Q���{��g<�ʝ
�k��A�>7��)QN�V&�ט��>�N���C%%�)sn��wk+|чK|�jٔ��f.�J[�ЎUe0��a�������>n�q"���pws�Py;vwE;<2�-��ϟ�^_�ȩv�F���e�O,�~�������#�ͲX(4*����k�"�@���������f7Ə�K %�G��jumF�/���3��/;s�Hŝ:N����|,�/��E�s���~�?�����ō���L�4l4���L�Vq��t%��P�q��W:`�x[q��.�&~dY��yՔϚ/IL��5��T�x �"}��/^�����.y�%�fZ�s\�Hp %�	�>,��Z�yk���ׅ��2�4ǡ�|�?"({>  +a�=q��H������P��zJCf"�nj[�5;�;?�J(�m��ƫS������?1�#�
�#����`��+��G~��5|!2����x�r��Tɱ��tƍ
\8���lw��R�͢���є���m��DVN
G�;�kg��q�	�s��\/E'�(�q�RΦ=��7Mr~]+G���?J[T%�7n��{��$�3e͐>�k�q����7��b�2����iW�]�(�⠳\�m" ɗ����߹�7Z���F� �+j�(l��c��j��L0Nxt�4�`��o4q�ڦ>�¬�q)l@D@�FqM�zA֚���(�\��eG:�{վ��30��Tx�{_p���wE���X�*(q�kW󽅳cU�r���ٿ�
Mʞ��*��	NF��`������F������dd���n����eP����w�S��߁@GQ��:UW�����������)	�Z���x5%bfG4�5A�!8CeN�~��?�z���υ궊2P��;F՛�7��vN�����<�����L��I[^q��tKATv{���'[�iF�i�,YF���`Sח�ɏv&���rOt�X?��aLa�t]*d�l0Zv�W��A�A�L�L�`��:ڤ(P��~nE�v��1;�&6���J��r"
�`n�T.�u�}�k&Ch>�*�k��e�U;+EqS�Ǐ".B��2?d !BN?�;V����2y���W���U��>���q6�qy�1���<�\�0�n�aLaWgv�q����9�����.}]!����\}r��)ͣ���=��j����R��	�V(=f<�k�fA�n��Ι.�U�D]^C$)$��o��{_MlL�dwJ8h���F�jia�mu�j���Z�2��>����F��^`�9rPӇ]����*�
�1]B�a�������Lj��f�:AI��ON$��6}m�&d��
�u�*s������cb� Qo�t�����R��$�f(��Aa���o�j�+M5�*�oh�U�g6��jk��qZM�?�f�O���M�������'�F�s�Y7͵�8�_����jܶ�V�G���ݡQ@����������h�6���>���6�={�u}2�2�K�U&�����bE��F2�%�.�-W�I�Y��dDK[�֭��1u��r�u��Q��և�||:c��/py䵚�ij��=���+�A���]'	��2��#�krX������e�_���-����u�,!m���(���(�����!R�aYki�kly�'ü}bT�������c��7u�'��D��	�ix%��+�Sk��&� )�f�&�*(&%�F?k^�HD&�Y3B�qtys �e1���|n����®�����o�1��+��;ٗjj�{X�c�⟏0\���)^�T�̗/� ����rW����Q�D�$�n����}���m����D֋��O���k������X6�����(g���<�����l�]?���4��O�X�k˶
��0����E��q������?Ǫ��C^L�엔����FU-H���y��thp�?9�W���.��B�>o�qb��������j@�f�p�]A�� DC�����`���x���ync�z6������y�4��_.ڔ���{6��a�8"Q�L��#��/#��Q�I`
��g/��������<q�I������������^�a7~f/�g<�Pƽh�=��-������T/&����u��z}�C��J��'��?�+���#��o�JT>e������m�R�r�[�}U]MU�i7���U떕d�&S�����C|���~�T�]Џ�?	���)�r�7�4x1��������~QD�yB��i3+�fd)��C�;�	�݀E��,i` �s���{i��7��?[je$<S���cY�`U�׿��*׿��c��9��*{�aV�.!0J�g#�L�V��c:�G�**\��(^o��(�հ�US�J��I� uoE>�	�F� ��f����ui�h���o�q"ZחE�h��ZK�΢+��&�������T�-⫔�1k�K��S������>��78�lvll��'�ITܔ�u���}���TK�fvl�HE@Q5��d	5
o�d����5�kQ�֔�Rq&`)��mT������ݗ��u��w�{��J�q�7R��A����X�7%�� Zz�������2��8o�ɻ�]C}j Ǌߋa�hqF%$$Ե�+<
����i_�wIGU�\�!^ғ�M�
{�~0��uB��඗+����T��a����$L/g�3�a��X��� FھokZ�N�n�K�A���$J�v\�n�l�� ��KGf����{��2=�S6t4���u��Ń6>܈2��t���~�<IBdtt��،ŏ%;$|����a��'#{k�@JW�C���غ��?  � �a�Aʹ�R�1YEPX �����K�6|��A�f�\�G��J�����:<�.@��-^KpY�%oou�]ng�&�����w'v�ݿ�'�U�ї�CA��?�[�/%��.�f��^amc߯�oŋ�ABT����15%_>2	�3��`�h\x������/��;^͓������ZJ=#��\��8NK��`oio�h�F��y�+�8Ō2{��"5Z_�(%������}�d�;H �ʞQj�M�;�4���n�Q_����a7��~��|�3��Ia���\���ݻ��Y~�^��✻��W�UWa�ə#�\�ee {zz�V�n�>����G�)����i6P��	@���T~m�BP���ؾ�u���2+`#n Aw{��;���ш_�$2�W��+��X��!毷V/��uK�*q��jެ��費-���.5Yc�0JF��-{1B�
��=|EIIY�o������@�:Y�U�<�Ƣ�m0�2����CL�Cp�mlR����>௦!<�����y�=+Ǵ�QE���zd�� c���:�=��9_�������G*�H}���q��������L]��͹���l�|���z�k��~\���¯�uݒ>׏�;��S������M��ׅۢj�ޔZ5kojU�Q#j����U�gѢZ��,�v��{� �.�D����}�?�~����9��s�9J=_
��q^q!Gf���*Z�_~��W)�CѺ_�-�&$$+�ᨊ�<��i.��8Ǵ�����xs����E{���G�Ը�{,�Խ6y�T�D�W7d圣KA�/���[Q�@��P!��b�Dv�|��~Eyu5"����ۯP��ײ��~����K���Ŵ����觸$6��½(�5��pu-Wп;0<� ap����ϧ��e�Lbu�v���ͺ���e���v���X�#pBh�zlNWق,����O�|�G8
�G�9����Rc7����X�4���uz��Qg��8L�:��*��N����p��PG껕�3Û?ĎX�i��f�"K?���m�J��cLzx}�t��G���2�q��L�-��7�_�PG�����x���0�~-,Th������\���SSs�{'`w����b��aT��b>J*����0g̕�>�es�zaR��#�t'a3�j��N$i���T�mG��>�l�yZ.�� $��z�*�����s�2A�#˕){�X��9]��͘��d�[OHO������AU\�ԁ�I�e�v�<$����2?�����9G�A���R�:��+-$�^�X��������7t��N�v�./���!gڰG_>��>RF\�}�.Q�u��Ӣ�><�&�����a4��f�����KV�l}�TCBҶ"�la�.(�nڤ��%+�n,�~{
[�=^7a)D��L���%?���;}�s���yHQ{E�D"7.��lc�T劌����=4�E4����ަ��>m�F $�n-P� ��c��!�b���r�������)�g��d��~�������踮gl�Z�"h�iQ'R�Iԭ�Z�
H
�g�	��ҥ������7���_�/E��͊��\Fl1%�O�Uf���gS6I��[CZ��}je9.�S�����J-�P��ƛ.�(:L;��E��J:����*�X��^��x�5���Zb�e`U2�l)���T�봸����c����O���/`�:�z�I��������c=B橨����(����g�Wxڟ�$�/H�gK���ݘ�Urjm�L���#gu
��m_��[?��|��[!hZ=NNi1zq��|X72����"y�*���K|��@\�t��?T1��	�s0ӝ���3��'f/2�}g�ZI��K�2�/C�V�"r���d���#l�d����P홍��Y��lgL	���ψI1t^��z]�^zeQ��,!�j����(�k�a�,V|��˨����Q]
� �N��C���*����S�D�����	���s�Z��}��ɟD)jG������S�&�}qs����y��3�
�.���'�A4h����`�j[�k����±`�E��M$�d.�R�����x��B랉S��Fe|+z�����lڂ:E�`�X �qa��g�&�/;���~"/Y����P��{�w�8��fk��yB^N�z����������u��Ie����^���D�����?��66��L�sb꭭n�c�ЪZ�oEd#8+��oڭ��;(��&H̀�;��O�T��
`Ig�2�#J����H��Z� ܰ��:��%������[��z��L|�#��ϫ�N���%D��{�y��jIF����1����oEzb#�l��:�6q���>\�_��`���ߋLD���nC��uk��0�O��.J|�U)J;#n��:��8Զs
���r'ӑ'�/{To�iڐ|���������!���xGT�秠��)~o�DV[���}W��߈�k���1�����sttD1���E^��3��X��y��X�=Lc{�K	��Cvs����#�輻�3;���j2�>k�����`|h���Y2s����KT��+��ȂuJ�4-�[��$Ҍ\j�r��O]�]d�w���!�XVyZlEf���'\��L=��;�q���.cOg���������Oš���.�-��̜-`�"�b�8b�C���q���C�4�B���8;Z���;��f�烼WG)�+�ߋ��L�o�� �<h�{�Iԅ
����cS'w°t�:�N�tu�@j����xsj^<R����D?��� ���W��Y�c����o�'u��
b:ְ���C����۫ߥ�)̷Ǳ)���ψ<�޼���WYƔG��C|��:/�|���U1��[�������8G�z�����o���F���C �J܍�]�
r����F�����k�>��
���'�*��-�J���\&���<��OM?,�38u�e��]E�z�o<j���q�<cˤ��<{Y�]��y���������
l�<���#z�̼b�.�*�x�p�����,�|rK:���:r��]2�+ɓ���K�|@@������S��X���co��j�9�.s��r�)�-�ފ�12������6�a�>������ǫ�v����^֓���K5KtV�������}�pY��?��	���_��y �w�ܤ��.4��{�Zyؔ��ύ0�+��	�<���jĥ42�X����8e�$��ڕ�n�?�l�-%[���֗��I���g.aN�C�_Z��J�Ը;�b1�x<�O�j�e������(�]~ki���WQRz��[�)`��q$S)k)d��|���!gD�0o<]�dwߒ����f���&иf�ēBpڂ�{d���o��U������"���=@�}	��T���=
�s�a0.�)���Ϭ�E(�CNc	�2�ٵ�}���?���:t�DəC����nm�K�<F���0�Y�$ä4��#W?	;H��T$&Yi�_`���'<k/ŗo
"�_0�x��@��<`Y�e/�7G�B��;�/�̷#F���j.Y2h�������6�W͏���ql�k�3�"ޚ��*�)n=�hf�����mI�}ڷ�I ��~���t��������O���������b>N6�֮Yhz�9��vY��9�"�6���7S�'���b�K��C��Ta��魍��=�q����J��h��A�?�5��X�z�,�BH/�^�qD���q�c������C�^�U��Wm���|]�4PGl �hF8����n耒}�i�Lo���G�=4�6ؘ��I��lnT��oG�d��4�oE|LA��Ӵ���.�i��2��(M���ֺGQ4��Ҡ(�eyRo~5a�?˿���0^��\n�+HJwW��_R�Z9`"2ob/���$y
9,�,2~��OnO�m�X��PY����7��Xg�RR7-�n5|���-��_hp�"Y.������L��IQ	()�?s$
M+iL.�_]@���Z�֬Q��u�>%.��4-]���&:(��T�6��T��xY='�S���OP���{�7�ǥ��vV����j8���97t/�hyς*��8��5�m�h�����E4��d���c��h�ѹV|*����G
�w!�$�͗�Õ�{���YX�Vp��&�
�pe-�PDs0p������O6cIp D�R.�(dN��i� ����J�����*S�����!-��䬸1�x�f$��@�mP�<j����%`%(e3}so���������d��<^[�S�N�q�(�:�`N�E�� /�T���/Q#�Fd��G��vա�_K!��T}i�bџ���������ة�y'�
�~r����d5�%��e��F|z^&u����Y����@�ި������YKk�i�6?͙q�x�]�/^S�`��0[
L�/�����* SS�¡�����%^՛6�\F����͗�1�CÂ�(ɦ������%���O�\0�v�A�R�����ӿtc�S1U��P�o���&�r��(PF��*>i�շ��!ۘO���+
�9��ח����
:$�mM�̡���_&��-$`R�f��k]7j_�\�5Ñ1�g������R��[	�gۥ�q	V��ϡYq�!H�9؟P%��2y�Y���~ȺY��OW�vX�xBG��|-T�tY�;���G�l�q��O$�թ��l���Ӝ�l��C{���'�ԢeK�9���f�
x��OAa��Ѝ���)�/X ���4�?H�eJ�r��������� b�#�9��A�[mW>w+1E��u��;��g^�
�q�\��{9����������|���M�' ƛ̈́�u��񞰣Q�^Y���c�b)�Dě�p��E�9ju�GsE�=�B�S~��Wى\�l������m�Հ�HG�In��,!k�f�b�#�v�cӒ}�� m��ju {Vw]z�/qu�NN��&����ZE��O�?���� v��-�k�mC|Y����[�G儙�e
m�f�+��� ��X�N�$������I^A�ӊ76JJX���'�������~�`��G|+�DC�8n��8����Ֆܦ�,N��秒��M�Mw�(�������=�3��-��g{���{��ʞ��bhʤFj�y����r4��obAhf���/��ux]��(�����<Js�]}�2�WQ2r���`#�a�HK���-�^�Z\dpԽS��k�?1�
2ϫ���lu���a���v	6#�C�{���3w֚�Tª�}�j��4�.E5�u��y^� ~FjlĎh�L��n�ΞI" ��,�^�ǥ�]n��d-6�F�~�$����xX�=�^e�dI![4k�3�&(#���πIv�8�Q��:�)->��T�-�Z�h�d{ZFq��T�M����J���je--"��Kk�OB%l����u�N��`�s�$��YKy���Jz��j�R�S�WU���TQ�)��9�S�ߊ��H�3�����f�P��IS~����"	��h��@�o�|�u�_کljj�h)`=�Y�w�}���^��|
 	�^�|G�ȍ}�݌��m�z��]>�D$�����\�СN�ͪ����'_�q�?y�vE䓁DV�6���K��vYHk�ݗl�"'��+	���hgE<%H�F��p�a��}/���ɷY��7��-���������V�����e�����w�{����������M/��?z���j�{;���¯K���&ce����[����s���)�+T��G5�� ռ/<�8���u�T�a�U���g��5=�zWQ��s��Z�9�XH���΃�z�\	�=�\q#��it�^��=a�H��_H�j�1���n�s��(�2��O���B��i3���iT$n��G��л�hʟ8Dl�l�sq/���.���t�U!}ι/.�M�|���2��L�R1���6$b]��vN��Aǅ��S|�4�� ���
�� �=���H���v���[���b̕���1����~^Q���N> p��F6!�x���җ�:�L�r��ԟGȽ�ԩ�R3�� �`��8 �0�nz��;��6@�Z)��NR�m;QNf��~,�ޖ��ھ�dY_x��B���sDD=��W�5�t��D`�u=��I���;_�E	�,���ܚHk�8���ӗ�/�4Z�ih���齌'G�.��PH-.���M~���]hl*z�_s�]kR����O�ݞ�>�L�#�I�k&�-+#b
�}�����Cٔp�5eZ?k����5�׆{��[C{���i-�ʶ���as׷���V����kYJBε(��g�J�DFPo  G/=<jꙋ[��=a�.!���H���;E+��=�WKL��٣����Bo���Vu"��nq)�4t,)L�#Q]W(��ks�8��Ӹ���z���i�2��&�4 �e�E"@�ϝ^T��y�#7���D�<;���ˮ�Q�`;���K�`3l�^��<��̉Y^�s�w���A��k��%_�=�a +��o��%<��Wh/���LE�����
>�o�xE{4�t'h��1/��Z����R!���LY�
<��_4&����2{O�y���x���+��Wl���G[�d����kA����$�]UX�+�%���^��H&��D_��E�Ć9��2�E��qHcu�]��xT�"hY�i���s�ՀvL�It����f`jʟ�r��5|�uN.[�����.!0���Gy�ܡ+вE���A�����;,�!�^�7e�b
yI0em�]5����qU���E/��Iy�R�t|�{̣A��pW8Q~tt� 3�{+!�T�0Ǚ-ݯ	W^�G���<�0\A1_���/��1��})��eNqFb��9���jo��
���p���#:oKO-}���>��76�-8G��͹� ������w�$�
by��L�]݆��g<M����A��o�4E�)S�q�&2bx9	�y����w���0&0�3`X�r�u���H�V L������U�֔�9��)$�6��qSKKIL ¯���C�ʵꯛ������� �@^Ycy^��9��F���Nq}@�_�ܹ,�	ڽ�x�����K}�r��;���qdFF�Ѽ�����( �*�aYZ�$�|�G���%��j����#��'�(�<�O������yq���N*�%hմ�[`�n�番���|�y����G��¡�ЕX�omr��������OH�=WH��v�d������aA��aQ<l�Op�N^zn����n<1����2�?.���|�!�C��N�gi.�m�XF2O�
���+��Z�xA/H��s��҇������v��Q�^��=�5���r�g;c�*���o�	���X����~+���P���C0�-x�@"�籶�͟WD�	^hu0�^w�kV�M*!0c@k� Z���������S�(�q9>�UͿg�Q��O�M��(��cm���.�wy������F5?��`���|�f� �,<�� 6՚:�=�'�2hn��'B��[9�$tRy�NW!��t���8�:�|B����` �^,Qߐ�;����ѣ�F����3��]��ʡ��C��D��c䈙�[�톿u��xA�#ALK�;��Ñu:�à\�Q�N�����j��U�P�g��a��;crON�d��K,+^�,���p�b����.n�z
f��I��E�y����a�U;8!�N�H�o9�����X��ёF�w1��Å^c�Pe�Cg��G���R�^�����n`�L{��!3Z��P����K��lT?HU��^Z-�Z�E(���wg�Y��@Ҝf+�����A���0OBQ�
`RI��2G�����n<��R��G[Ӵ��6��>�c���
3���R)�%�
��C��J݇�R�3����'o\S����0�-?:fw{�q�ס6s�ς[A�,~�K�����NN�!鎓7�L=p�4�"Z�j�A&�˟A�/���fW1�4�v�O��]�d�<���ݧ���xm:���9��^o~�X����*l����,K��v�z�`4������H�j_��`��\����#���m��Z����r����@�,[�PD�S������G�O�/�.+�䀤{��@�j�^�iW�N��n�MY�UN�Eƣ��'����|�m;9�A�c���q��d�ۆ������^mx�V���4b��'��O/��O<�������x��<�n>�]t�L���<�Z��G��-��j���S��_m�x����W�^��E�t<�'���ł4Bz�z�-Ɗ���~Pы��}�P�!1sO��-h����վ�WA����wz�xk9ˋ5����-��
��=���2#�r:�H� ��C�SȎΘ]w��c�$�T�����-����2b�#�O�_I�d�Ҡ,�O0Ζ��;/סLb�ō~���~Do7��x�R�ٸ4	�ͩ�0	И�!k/xD�Rb{��Ίm 3U�E>۶H5�Gm~����9@i��G���� u�͋�� �����侂
�_ BA��ohƜ��.�9P�v���B���a!���h��E4-w<	6�����F�V/�r:�?{x�Z>�a�t4��Bs�c�%e�*ww}����y�*>�C���YsJ��?�\9�5��"���ʺ���姀�]���7T��w���?�s��`2���U���V7Hhf��<�VΘ�:�����!�n:��^��n�Np��9c.���Ϸ1 �2�X0�7�7�Ь�XJ�}�Q�Y5�χ��[�T�jܥ����U����_�ks��k�?C��pDGWF�5�T�*���[�!eF�0T��{����� L�����ހHDkd��u�s���s�o�PbQ%C�2�}��O�����/��,.XHc�+��������_�p�z����70rR>�W��I��p��p�/�C�3ه�)2Qv�f~�9�ɭ��#���83�2�
��3~��D/N�*s��e
�����a�/h��@T���mg���wڄ%X߹������(@��L��`�5B�z�%	���KG�E�|�$q[F,vZFCdF&H����l߅ �;7=�l�\/T ��PЎQ	�{m��@JV�w��"G�p�ۮ��]Z��j|�W��ъ'��m (��]�G;H��2����D$hj�>����Eܗ=����+�/L<f�ct��T�D�GlW�ѕA����ס���Ն��!��E�&_lKF�u|G��8j�|˖X�Zt��&yGE�Q�G���yB�n���l�@�nބ��O�[v�hP+�E��)�I�D���a�g譂G�=S�xE�}�&�H3��J%�O��*���]��\k�Y�o��6np&͟@�\?*L�&�)8���E�RG����a�2X�>/(��2:�	)��|G>o3;	z���8�KlvF?�A�T�k���/���jI܏�]���x��p�׼Z3����U��<�M|#�~�mV�.��	{`�쮊�iӇh!K9�����y�X���%�Ϛ��+�1g�5!%2�,S��s�Kd�_c_��>OHK�:6����`v����|�h�F�e}�����}�횙88�"q����zw���Gd����g��	!�p�"��w��"��@k�(��p�m�=::�=j�'"�^�M<M��\\�����&i�"v�K�̌g�`x6��l���*+2+ƾ�͘ʵ����l���^W[݈/#+z^��dN*�/�1.�M����?(����l��DD�i9��I��j~r��.D���!n�#�N>�����P�o�nTC�n��1�k���WPU�OI�z��x�F����U/�c��/��	<ÍT��ւN`��{���2�=_�������^���<(G缈s\.wN�zw����L/5�i��5:����V/dΙ(�ƈXo?�1q�o�=;�����6��=���j��������r[',���-�c��'w��9��_05
m4�'�D�է��6��6v�U:�!���K��Пջ
*[��q,�3��0��*D�q~����V�QU`� ��\z5sD�0i���t�ș��������M��uj<d�Z�d���]rL>>�:j���0��(V�/,��ܥJ�yc#BM*�MA�#'��+�;0�6���[��l$`u1Jdz��2���d'��T����3��~�3�9Ӻ�޲M{��;y������:�C��%����6y0US�H}P��9S����m�����������L��c�贛���n�r��~�j���u7d_(�Τuq8R�c�[J7�#����+0���S�K�ĒtG��@7��K;k��Θ�Kjxc2�sQ�^=^3��q �4���e�-�>����/{�<��H��<�؊��q<Czg�H��9�2?��m�E#�R)�V=qN����T�4#���|�m�M���2�׳f��u�Xr�ַ�F��Q�Ƥٺ%�?^N���[�鄓�^��"�w��^���{R��P�mi?b���"f��+W,TR�M�-Iyko��#8�q�ܓ�{X,�g2�cE�O��ԥ�����hl�,$���*8l�[����~�B+��h�����ᖖh�#�Ass��Åjd9Z���\�VyTN����Ok$�ǎ�?��hd@��6�c%��%�K��cKS4g��M���_��x�AM�������y%%U
o��~yw����'בy���p�jF�����-b����毗=1��%ԟ��4�k����sJg�X��i������ͷ��@\���e�����Eh{(��/�X�9%�#a�a��i5Aɗ{.�M[���U����4���gB�O>[	�t���\�
�4��r ԑb}ހd��o�2����g�Ś�u1��ؗ��$B̜WI��.��
�u�2�<��E�tw�������XonX���Pe��a?vB��k��2����\��ꡃѪ]���<-�6]�8e߿�-ʺ	6&N�[��q
ۃS�b 鋅~K��bޢ�=�> �ݵ�Z���~JD�KjjAG��{��6�|�d�i�*p{���g��
h�E�_�a頬�/�2�(vl��������߾��X�:�W�r���ү�^k)���H(��bu��k��5je�Z�\e�zsX�,e�O�nѣz�}dݼ����4�1|��t�ǩ��~B�&u|���/��_��J��,��~W�6�՘�M	*TP�W��Hw~��%T�FDw�#gt�� =F�כ*�>��2�l�_o�F� ���~��ʏX���w�I�����SA�
���u\�����}��hB���˶�sh/�	������kF,CpT���9���xB��� e��X-��r3�go*z�nN�Kq�)�ѧ�}� �?Oܳ�Nu�`d����u��J?��!�eaz=VnPQ0(������i7?@�!���%noJ�܌��e�yk(:��`\���9�d���r��-�����i�.eޘ���	THS��qx�kX�����2�im$�LƦLý!��ݙ
hm4�G�r�X�>��TJ�k�.�l^���D������Q�2W����nN1�wj��ё�]�>2-^1|�l��W���$Z��6RP�8戮��Y�
��2���Zǉ_�I��8�b�s�|�yj�~.�	<wH�SڱϞxd_�9we�A�9@�9�$찑�ʤ ~uA�:��V�����.[��Ꞔ������Q�4u���gXt��`�uE�|�v�sy�>��l��NNaBT9훾Xf]j�h���dߛ�J�%W�LoYq�QL��6����M��V��7��O/܇�R�9�6�B��#�)`ErL~B�ґ^8rێ:�̿e�5���Gͤ��u�h�*.�6
y�V_t�P�TG��Y73w�����hM5���2|H��$�Q��W 56���t��ڀ�jȔ�,RY�J_q�����1�즿�����l�ighZ��H139�`�����ԈVQ'SYq�h��5Nn����k���e��Aj��ҳ���)�����p���[Z_��p:��Sų�a?�w�@!xѯ�~x@�xA'vw[��f}�Z�W��6�2��=��5*����TIpn/��_8I���ZI��LiPJ[y-�����x��|W��\���\�H|�KD�9��yc�+g�t�� J��Zv�V؆qW��y����-�{N��5���B����N�{Y����a��>��=�����l�^�R�� WS�����Z��a'�"Y�U�����Un"G����5V(\��0*"��{h���[�^�ֳ`ꜫ��'S�/PCy)<W�9�O��
��p���!z �8<�A.�q%>�D	2U�H�{_/ �������1��uU|7�H���W������][CD��������_X�~ӽ(���VL���hڹo;��t��%bs��ْɚ/��{�8��?�y�׷��2=�`��r����, ���M�'R姹�;����O*�2�K�5�����T����bSM����o#��[5����3qɌΉ��j�-�-�9��ֹ9P�Ef�BMҧ5�����hfJ�?&�p��ï0j@_�&�=�˺z�\	�U�����i�b���)=͍��<�a����ӆ�&fyw��<�������:�j[�8��%
�W�aJi�}�]W"S�/�#I{�1�w
���H��i�#X�36(Q��5�g��;��MS��S�.��[�i��^�17>�*�W�q�pz��'���2����O�J��򴴟��9���߯��W��1Rp�_~�e��Y�/����b�/UUq�<V[r��~�J�]|�A�7�����r��s��x��w W2v�N�OZ�������"H�#c��9^����'ph{��`�u�2pk��s����v��*[L�|h����C?��S�.��
���Jf�L����L�w����1��_�\e�t���Y�XU&�pkA�O��;))8��)(i�LBg>ǟ��*v(CE�Ӈ�P%��i�F��⁁�v0Bvyy��� V(/"@���v6����q��;"3�J椗�F>,�M�SغQ�c��3�dӈ��a��9��x�}!�0�镣��C�"9%/L�n@�+�!Z�s�È�Ǿĭ4n�}R�c���Q��ĥ���ޗp�R���Αډ��J����X�P�N
��B������m��<�>��:ZZDttt2}ԟ��nz�2��Ne�|��'Wn$�%�勑%'ߋȫvg��,c�'�!�n:�,^���X����r�)�I(,q����b꩏ÞT���������[_)"�":ucߣP��E����B�دǐ�6G��ˇ��N-�l�*�I�E8;;OJ�S��8����������y�?�����)�Y02�P�]�
�����u���1B^��m��}��k�NWz.E�:j�~m��@^>+s[uS�oii���D�z��p�̈V��r��VY������w6��i-:F.�"���@ծ04��!�@e�W��%������*��6��M����3�?���~�z��rC�|�<zws˖.���N�]�}$���X�sCt@�n�@�y��� �����ku���_��]q@�E����!Q��6�k��s¤|�B�*y����~^�R�'�/OmΘK���
u��*�z�I��J��r���F#���>K�|8�b�/�����f�����C>~�dSW�8�ع���N������5�9�:j�_L�l6��RB����k,������[�x͚ۏ��`��9\'ؿ�jT@���ԴM�D�rʄ����^��mM�\�VL�w˖:�59s�'�C,���U\��7�?������ZX��\(��{b�DYT	�^�6��5�=���Xu,���%�ԉ�2)(������ɥ��*�i\4df���'��<<�(4$y,E	O��Ж�@�7A����z>���M��ү�*ӷ�aG31o��z����� �u>P�gh�0A)?�P��<:�'.���'��˻_�vf�� MG?`r�%�ٲ�ܔ�ebL���I�rJz����!�g�_$}M�s$� S�:�u>3��ψ	���<�qo���+�5m��4�{c$,��861��|���)򠸵�g���p����C���Tܾ"��1Q�J��B݋���R�+��װ��C<?�_C� 3���%���է�:�v��I��ݻ��0&���R)_����@�I~3�pN�r��2�n��Q����VR�#B,2�������WZ:M`���g�+j�NtT���p�3??����ۿ�Y�Ͳ�S������(�Rso�h�2��}��x���\��B�%���~�o8ѿ�s�F�o�o0p�8��DP�K�;'ocJ��lҶD�p#à1ݱ����s����5��\tt0a2�hȄ�8��y���eT2�,����A�P.�C8�I&J����j9:j�{�@g[8�����Wg�a��֛@-"gg��.�T��H��a��s�h����,+�,w=i��>��v����� �`�w��{aCn�|�>��!X$��j�R�^_�e~inn>�f?�0�=�Z1���$�[ɸh[6
��jP��@�����S4��):^,��5������T�[�(8f�:&�4:o��ɜ�G�������8��l���������\�j������󆝰�A�L�?U'bu�!�>��H���)-�7J^mo�S�0�n;��8����F������׏�������3���S@�����HS����b���2�r'�V���69�����ʯ����խ��4��,�lI��0�q;����e��,#��v��z�ؚ���U=���VH�1��>�JBӨ�E9"�1���O�1uj��ɛ�^��ĉn:� `v�|di���(|�������'_�o͔� �T�|e�@{�LY)oI=����B͹NN�u���ޒ�������4��w<���������������2�@�I�+!T�������C�w���=���ze�h2#�X��,�F�݅�-���Q�.��D��H�ׯ7��m���7�/��eS�L�,����]��/(��� �|�|�E���+�w�J��������v������P�<���_�]�~�/��s��5��x�7m:i�P�P��\Z~s`�#`��F�N6��c9<�nn0�%�ܑ?�{ak��Q{��_�*:�9���m�X4$e̚�H5��fHf��g�ΘŲ`�U�-�.`�!�v�ɓ�Ց=�����������޵���AB��E������������_�ޟll���)jhh,,����bL�b�X�:����8�u���@�^�e>�-sj_�g�.��cR��:���Z_?��,i|Y:{��?�������6��6~�`P�7W'j��hGZ��
�����;ao����B�_bW�����������v+���������k�p�,fo&��aї9�����%. ?����c[�-m��Fc�;��_�[މ��X;�R�����"�R�~���K���������}mov��v`s�@�J��9��oo��.����9��ʜ�>�"u�B���+�J6!u�+�w+����W�Sȷp>�<�JP��x
[��;�jK���Z���2(���}�$V��S���)��f~��^�n����ɸ���3�=��bQ�^��>�qb�� �bjF۫P D�k�6��kZ�<
ٕ.D�5cvC=�����d�/"�}Y�����[Qɔ8͆88�r�XI���U|&�2�1,�RP�����
�>��i>�#E.��؀���z�ʧM�U�~.��K;)RJ���1����b�ڏ,���qνec\�c���n���P3&�1�Ҝ���\�2�j�%pJb_�u�{M@�ʔ*�������4Y=�<�?��4���y	b��5�������H�<�p�|H�s�|��v��D�wvt��� �j�ϴ�f�� ?�_ҲI`��U,q����﬌R�UN����?�o�s�|"T�C�i�\Y�w	��V�81�n&Bٔ2��5�6��	R��9��Ÿ@����`��G��5��ŵ1`#�d��h�K{Z�fA����V�Dr`ܙ��c�T����OJc����a4�Xm�fƽ�r9��y�*>́+����g�&�g�uǳ���#+i&&YǃqcUs�@��S�\�"U�s���7���&[r�o���@� � p�2�/�ӛZ��������h��/�"��վ�M�ٍ�@�r0y|D�۽r[2Lv-rQP��#G.YQ�������ߺ� "�s���o5c6��~�"A�O��Ȧ�qQ�������tqU�_SJg���PsF]C��I>�k=�2L�D��0��K�'�b+3׃�\�nT������P��-n�7�b����E"[�(2�Rc�K/w�?K���c8L��@�����}4�8�e����3Hz}�+�֭!�� ��Ds�����©;z;��SĠ(f�`�]+WlƎ��H��G0�
T;Rm�hr� �g薉d����0����K0�蘧�$J�:�@4o�bnC��?K0U�FoV���M��@����~�9#M�?��̄Eβ����'|l��M����	w�9����{� ̰���OJN�����$1]�THg�)U
�?7�6p;W6�F����`�+b�g�r�ǭ-aeUȏ����KWg�!Xh*�fy+�&���|���{3ڹ�zΥ�*B6����4*ս���k��'����	�˅��/�BeN�fҿ�ɣ�3�4H�D�Y�| u����$M� �������wk��]����$G`g�����0�(F��Px��p���@n�>TaÖ3�P/��ɡ�d�^���6�����_ƕ�_y���G�3��� r�C��,|ϛ��w	��b8YI�Z
$"Q��'^7�X�s��Cy�	.�,��)ۭ�m�Y�$ޤ���'�(��]v��=��\��?�x�h���b�osSKwR�[z��$�������������Q]��sZ�^�E&�<��=c3E���ʟ�&��~��o+�ZZ�39�[�6r
�tDD�>���oֵvE:�y+bf5����}^}�a������/7g9�ƕA��n|O�|90����r3ʈ"��ϝ�CP�՘��q�3��w�y�F�՗�x9M?��v�6H�O��N���Z^�Ϙ0��*+%�Z�`*��K���P<�C�:�7.�;��lĤ�Y�Om��1�O���ED0�N{=�m,��u��k�7�ρ;��__���
p�#!�t�����Q#�2㖘�C��"{����_���JO�u{�9x�ɤ�a�����W ��5����Cp�Cp������ݗ���K�]���	�o7��^=��������眾�}�)���<-V���C�p�R�0��`3����g@��g�,"��/�H8�����$�J������(���He�Y�nv�"\�8e��,{e�5d{����7�I���
4�n��@�����Z���w�sҺ���_�؄���I�һa��I���5�l@:������?�6����I6�߄O�����.R���7��fbS~-�f`C���do����k%t�DR�0y�f�r���@\H}�N�KB|�rv`n3N.)��gf�q�˰S"�;��?�.Z���#��r?gB��:�.��_���w~�*!Ŗ+^r���l4B�{��0�Q�Bݞ�Ľ��m����gƯ��b��w�|̇3W�Rm�9n�lW>�F�!*�w�&~��}�ڨX����f� ���h�q��?T`�LOǇ�e<[����o7�LW.�����������nñ�*lL�Ӳ�˽��Ł�/	�p6��p`��z&�7����y��k	�E� �A�<�FƟ$�Hї ��(��+��B��B{�!�ş�33A�ӵN/���)���%Z9 � �5���iݘ����R��kU��I!��Uӳ 27-Y�����5��KO���ޚ��\�UV���׋�#�3����J<��3w��Y�+2p�#��%Pr�5�چ!��vKO|�8��֧�6l�;�ZlF�Tr���fI�	[�B&g��!^FW{��d��罐R\s@噬C��뗆Dga�:I)�,j��)	��;'������rw~��+d��g:�(�1�����7l�|?���jo����cc�ǹ/�J����r=�w5�%�N�DW�nȺ�������PY�7(7SGkʡ�l�c���K	a;�!�`S1hw��m�*c�0ºI�J:\i�u$g�x�E�Z� �r2�#^]HwUgQ|:���!e�Z�p�3��q`Rc
�3pV���)^X�рb����f��?f
z���ڎ�5��w��*����8q��u���m��Ib$�niiD; p�]՗���|t� Ff[-ߖ�lX��4����?���CY['���>:��ӵa�@Q�_.�35y���B���g�L�(log���oJ��{�w̨w�$*��ʐ�n�PW4)IV�f�V����_'w[�����m,��V�>�p�l����D���J:R���W���7�B<$v�/b;�>���~���Х}��W���o#���5j�/��N��Q�2\�`Zx�����r �'Ț��AN)4> S۰����YfYa��MRc��t�ZbTV�S�}�h}�a(�e�~ȡ���)����ř?�CU��!a�8��H�,�]��2�֨�����qa�9���K2�D�m�:�t/R3ݛe����"��:m`����
��_-�g���Y$�����Α��bv��R7;>uc��� �7@����U\k�>��ў8���Z�;ߴIh�r�%���A������-?L���;j,/,�V�E�'��ӕܨ2=~��h'+��g�Nl�?l��>�7�ܱ��W�P�DCC��;B�<��r�����4��hDJ���>1_~�5hM�]k`-H�m�΁�	��VS��cI(���	�� ��I�f��W^���)��G�_J���g�ڽy|������� t�z"I���{�����p�����I��t%D+���ҡ����O�}�7�o8���A#iK�6�C���*�\��&���吖����Ď$�����OeC�O���|au��sc�\)�a,OGL����m4_W	9�,�ޥQ����Bj�r}��e�"Q��;(��o-���|+��Z�c�����%��O��YX�Z|?97X�t�a�}�>1u���R�xk~�4�ޔ��)t`�Y}JCy���X4#�k���i��_�Y��0R��e�״�4��Z�!J$/���6�L+��n�:�o6 VB��!�(J�P�Ł��)ѿ�:��ąg�`���Q�"�0��G+Ni�h�zl�S�!�%Ov���5,��ŊC��P*��uo��]�<���!�Ǘ8�V�����6#��]]K����c ���Ku�^�'��ٙ�n������^�R�ꏇ���3�%��E�tv�B�Yr>��Q�Br��
x�`��9ܪd=��JTdHj�/��c�������v��t�P��ׁ�u�۱���!o��eN��--5��V�[zMw��QS����K�w,���I�O�IO��_�W1XN�K��t�^�U�Ώֽ���*�]������L����b#c�����v�fyb��ٟ�2�:�4���f����X�=Z�������@
�,������(#�]��c�^`�zR��`����7���QL8�U\PŷN��!n���O*��Y�>�}H��z�I*��=< �����-?k��$��x�/����]���O���s6�J���L?E���8��
���? ����wƺ�cO�5��gLNB0��,(���	�ׯJ9H'�i�w��0�#�>.�#�%Hn�n����|Oօ����#��啿�/�����~�k�X�>����z�����h�<:r5��ǩ����~�h���+N��+��ǘ�!�qcI�:܉䤏�a�4	����V�4c���C�;�G����y�!���X��y��{g��<���|k�U����A���,����ȞVD��s#��A~�,������>�j/�\��Y���2��OtG�ዧ&�>Gse�{Y�NGe?��e���@	�����Uu���i�LF��v�9.�B +sVY�lR䉅N9����h�!�G?�7H�P�=L8:Y>�^-�ZW�,v��е�8S�I����깛��[�����'Bt���Fi4��כ�U92���f���Rdu�7@!Ô\ta�?�q��G��w8��<9I8ć�ꑰ�l?:IB
�=��΂QX��0�����N)t�����j����27R�-͛0�I�c��;�M����,���s�#y#�R�.�C��&��r����&������c�?]����mѽ&twE)Z�"�(�g�9mCT4P`^��h�5�/����ZM�Z��-��E?'Ӥ�^��%��dt�M��N(�|i�q&=�i�$V�fd8����_��:]�ȉ�},!��hf0Q�	�|/��S�w�ǡ%m� �@	���qxtr�ޝs�J �+Bvu�rc�*����q��[c���6$��EMY���@0�����0����/w[j�y!j�|d�r�2∌�Ƅ��F"K�DQ��_��+S����V�pF\A`��	���D���ջI�T������<`s�ͷ3�B$��w�:*#��O[҉/>�ŪYf)`֏�j�\�T~�1QQ�G�����f��o/�W��+
�p>��[��m�<k����x�L� ���)��␠�^e��C�V�u?��\�k�D��t�pe+�\�����*y0�W�c��3�������"���i�d�R�~�������+�1!ŗ�grY�K�:�BU�Q�Ws��2��G4c�N~S�L5��[��($���+��N��Q��R���m ��x��f/s�;�O\<���h���n����#��� ?���eտ�`�JPs��ԗ�tp~X?�ܰ��,c0��K0��!�� zˀK]��+JĎW�|�b�ss�2o 2ڧ/C^�](.]��Ѭ޹ɢ��ӂW���u�0=��l[��Og��wv^�8���`�Qv�؟���\`��UCzP�Ҍ��r���r�#�k��H3���9����2E��'~k�@W%�SLS�}ZᦑV"`��6ZS�u!��ߠ��*�f=�������~'�
�A�@)�k�F�}��k�{���؋f�}�H^~v��U$�ѺN��D#[A5��5�Q3��C��q��wgt�v��o9u��>��=-E�/Hg9�u���.�bش�fE.�K�!��ŀ|8-b�7�X�9�j}�˖�������"���*�EG�؅�������2L���ˆ���߆"U?�%�����ᬥ4�Q��/��rPR�qq1-�W��I�y��TxY�p�����6⚧#���l�k?��T|�nk����P`�]D�2u{���Y8D�d+a�i&k���F3D��T��'����	��.w���FB0gJ���j�
��2��.��*E��G�\��(o4�*U�z^o�>�Q�����
����O��K��6}�ڳ��9�Dl� �2��󅩹U���0½�4�Vces�5NgY����T�Z�ttML51%\�Q�nRe�KXbᛤD��x�s��'��q7G�,���t��3�ճ� ɋ�=��PB̩Z��Ω]��=՝|��ԭ��T�������Iq���!4ԙ��2d�0c�-'H�w_�M��Kc�wsh��cZA�E3(
�J�)�0J�h}����5�`#8ӑ�M��"�^�|����t�x�ǋ}��b��Qk_?������055�}��}���=��^)��y~�1�jYQ��U�P�r{����KKu:]%>���n"S��ݤ�HN�-|����1ٟB�����ܵ	��gXHG���i�|�<4
�~��u��iA�o׿�2�#���ޞDy)��t���Y��!���62D��?l��o��)�� �Ռl�ܔ�Z9!s �qZY܉�V�|��eL�u���EIw�v���姵�m���� �F�-���X`�ky��+��]UK�_��/} ����o��/��8�gEo�'�vP8��sGt�!�?�I٭^�?>!w�co�ih\v�.������9�����$��#��f�Њ�0 ��%�1'a+�*��]��"��W
����IyM]�I	9���c^�y����EE�J���������33"������~��@R,�,�۝��`��U�jD懗�h֘��9�v(�Ҽ}#?
Ӽ��#�7Uţۥq���z1�5��ֶ|��o@�	���X�ZZF���I�Y�Ʈa3ӈ�غ��o�#� �����J���n|K�O���?m/�X�����y�|��s?�x���;�aҌ8��d�S�ݭ>��Jt���,F8%p�
��=ɟK�aխ�Z����jT��`�n��r�pn��/�κG�΋���qޅ�г���3eBV,��ֻ� ѺWɝ������0c���3�����ď3|���鯛�v�W���Ъ���GCN<X���k��{q�##�4;������}�e9@T-SGI��;��?�V�Q�|���|��og�G �Q����ew���~�=/���X�hx�o�O�lT��N��ۅB��`fј�0��Pղ�Y�=�Z����^9C��t�LߙZA+
k+Ԥ��`�yY�B��[��-.<+`��D>l�e��N�<Rl7ٴ$7�<[�"�O���t�Djc)`$/�'���4I!�%,>~]�Ce;���6�QU���(X��(7��T�\!N`�U_~Q��������3c��W9��!��6���*fI�4�7�>��n��X�����>.�:|��)��������.��W���.n�w�z�|\���`�i
�|ҫ�dA�����0t	^$���_N��l�d����@^ir<�װS�E�(��4�4��9�w����s�_��:(��b"
b6/�_uUF�^\z�珮���[���A��]b	gH�.4}po��ܪ���n�}�k��m������0�5�����s"�:=�N1�6,�Ҿ�`�v�g4�y��yl�N����_!�,�s
���3͖��S�	X�۳�����5�����ι�uo��[���ƥ�՜[�Nn2��.����EV��_��C9�Ɨ��H�D�Z�LL�'o�d��nd��O�_p�w��bS�r��}R�4�7FE�e�{��Sb��ik��6�\k�.��*oC�������
�&�g��������.���N"6�G߃��jy��qk
-��fw�?(��P�� 0(�u5�k��iw�,��D�꯰Q��5<e��I,�Y��6��<z�@�A�LUM-��j{�đņ��൘e�Q^�</��\2�a-E�a_
u�&��0�B_ߏ�@x	*���3ysSy,	#RM����/�`���BKl��+\�t��
��{1�&5[$�z��ye�l�:]���2�vp$�Q�O��0�}��'��б���6Gǽ���~���ʇ����qM�o>P��F-!p�Y�W�H��`�n��'����ΐ�1���6����A0�~�H�I!N�uҨ����
�YQ�򡘜V++���UV�k��շ
�&+����� ��$�[������&��(X���U���Eu��B�IL�O�d���j�PC\XQ�j�I9|��&�l�*L��Z���n��ZN�j������
�rՖ+iH���w�6Y�a��ly�ȹr��A�8*����]���E��h:��K�H$����u��Ch���(-�]��R������D�N:��*QN��s)Rݻ���%�l(x�ߟ)��wvB��A?c�2d�do��u�::��qs�0����Ǭ�~����&�Ƅ�3�n���[0�^�:�_�IN�X/aw���y�#���Wn����f�S.�Jެ�'5�������\f���wG�'��y��q�X��oOM���Q�����,�����N=pE�Br�~�n
]b>b8�i����s~糷G�'o��b��o���^��Ja�&Y�=�k]^̾�{�@�("'��˭z"ڭ��ߚH�Ρ��ɥ�sQV�i�����q'��}�$��[���ף���TD���c�z���}p7�Y4 {BԜ��o�v��~���g�����VJ��W%��jߠg\e�Mx��)�����"�RA��< m���@J�f�A��h ��W�ZXV��(�"|F��F��B�H�9r-AD��
꓁A� �����R�>�vb ��b�(j-=����޴���}yFp��N��d��s��M[%v�ַ72DjPbON��)k�DT����,E�H��=�8^�t���?�R��� eQ.��/�eN��N"f�����2��+���E1��#���'�H轤ω,�*uJ��Y�*b��p��vu�3���Y��Gfꉽw���n�0�[#�8'vs�����}�ý�H�` ��m
l�:�S�W�.o�	ѷg"c^��4�H�D�T�d��ѕ��$��ͷ$��H;�A��������M8�4zH�K��g�m��1 _�u�{�)y$ǜP��q(k�5����l#�V����y����H�́1����V�����@��@�|�&��m�w� �����6�;��m2[0���B�5@nln&~�Ɣt!=:�-�`M�H5��16���ףF�2����]#�hƑ�iu����588���XJ�WN�w�gνʉe{���E���@ �9
�&�\MC	����PCn��r��J�j�B��j���zL�����[�(Ur���)3Wp��R���u;>Q&c(U�(�w�.F"(�{
��.SSTt�9��������^�e��P�O��Ӹs������ޞI<��#B���QZH*�j����$�
8�,öe#L�R�9�%KKP��	|?rJ̈� '�ٮxgN~��p�]�X|O\e�ǹ�p}�j�W�}���:T�QZ�%��uQ�}�(��!-Qq{/����eMǰ&�z�-]�e������8�X�ˌ�|��`�<��(�jf���^$i��#!�����Ʀ7��^�ˮ)���e�:��bBPwwt�	��7�Qv����*0��"0n�&#(L����N1]CbL����bTV�}�f�I0�}�R�0�3܊�P~�EG%��R�:x$UT�G+��ܞ�ɪ%�l�i'X���U+�,�21�Ƒw�ߖ�T�X��L��3��%I���aq�"Վ��UR������͐>:��:�t1��~���k<l�&��.h.0h��,i~��#��N�4�Ir�ΖZy�671J��A6j����H���n�4���և��}���Yjp0t�^:�i�K��&��L㧬��i���Ox̪Rh�Q �.�.|6(> W�p��hG���=C��#����@mx�5'I��>ё���9�a����ݟz���q����Y@$��p����چԣ$5��1�z�z�}#n>��i�@UC&W�RQJ`� ��#�E8�����&!���	��������	�.Q�qr
�z�{�������L7�}�?�ǂ�@@�9X
�����s�h��JgՏV��X�����M�'�#�'�9{��ju֚C�!I,,[�{s2P������Ć�U�X�̉��+���
���Oϕ/wRP�����Q�_��*8S�BS�U��b���P86��� w���$��'Ȍ{�c7����⪨XQHu��7�o����C,������J8�ǔ��?���VG5ے����0�LM���}D�?#R[k�A�'�-ނ��E�����G��72ӥQ�̇�?���Jl
cj�i�ƨ��m=����8�q��@'�[���~v��	6��n����C��p���$�ؔ��|���ӣ�����] -��ڊĞ;ؖ��l���.�HtCҸ<R�4Wa=4@*_P��Fm�Q��v&��SK�I$�zg�P^�n"����m��r <�h�"v���/�`KwBũ�ՌTfw-��wҊ)�~�߼��W+���$�+cq��ޑ|������;~����g�{��}]3۬�#h�'��w��s{���)�����8 #�R�
�t�WW��vQ9�x�¤)`��$v�mL8�{g�$![��{� X墲)�QTS�9�~��צ�`����T�lgDϏ���AF�0��
ط���k��c6�{���`�����������/���.|9J�4�r���Fb�I�Me�%:���0����r#�])��������F�{V�����âGӭ�5�V��;hk9Y��hnۦ��E��!�g�,��>�o�2��Fʯ�G�>k�:�t��Nnմ�L�[P�]��3ɸ���a�p��߮Tօ�$�q� ճh?��+i8ڟ(����$PL��G�_{�^�i2~���(��G��Hw1��S��ف�M��6�G$T����b��#$ 0�n>�+͒Z�c�:aݺߚZ�+�{�(D�u��|U��YF$HO��TEQGR�.kE*�+n�f
ڟ�t�;]��h���,ڡG!�3�\�.����dn���;�<�֫	�:�'��}q��߼<a	�Ka AQq}5|�&ܰ)M��H��DݻS[A� �:���Y塕&�/���̀�o�������?�Z#�W�ۍ���|�����eO���?�$r�M:m���"R[;I���0Y�\�B'��$9Am"Q�m�'h",fԥLA�:��D�δ
e�/��� ٌ���.g;�T�q%W�OU'�O}�8��.�c�yn�����/�13y6B��CU�Xi5��#m ^�@� ��㶄����O(����J|�iWL�c�ۦ������������p����w��Nz���1�K�����E=��}jJ�ǳI+�f�P=F��ix{j�n��
��*��~V�KFІ���Z��뿺�c 7����^"(y�0�r}g�UGz`�����Nvu%�x.��a�����p{���6�>8:2>�~����8n԰��ķ�����g�5��! p���������v��Sk�z�/_AӦ�(znQ�� ��t,؄Mx�ݧV]��p��K����p�_��qҍUT�7��Fj��0XF7 lߓo]��r(�3Y_ޝ¹�n�l�(�o��چ��]�@�2Z���({rf`�2ع�[^|�'����O�וE�a7�c�K��k���@NzX�6Y��9_Z��!ߛ�:�ڙ��W�hy�$Í�y<�5������Q,������k�H��}I����DD��b������k�u�'_%$�S��P-!�G�] �WJ��~I�c�/���1=T�C���8�J�s�dℭԞҠ�v,W��<����Ϫ��e�����w���:��ᄢM�˗����s�rKI��C��Q����'	C�C�s[Z��AUϡp�Sx�S��Vh���!�.�:΃��:���-�8+�o����#�Je|�P���dl��ZH��m��� 3/�0�����m͏��y`�G�`�iz�!�KA����P�����<��"qC
��q�تP�6�'�8O.6+�t����]S��UI��XX�Γ�ڛLd.,'
j�j���E�R�t|���xN��kB7Fq������MQJ���dI�Cgc����~��k����o[5���AA��sZ�u��)���O�9�$J��P���A;��1��Tp��B&���0ݳݤ4��"�k��2�+(�&�2��Pc=�����A�	�wn������F�U��O���.YƳi��#�r(��/j�o/��r�6Y}6�Iμ�	�n����a�U�Sл��B��╨�&:�`�	 ��<kF�?ooo� (��d�J�<�lo`B�6���󆤽����g��"4<>ٰ���7���B�ͯ�v_�[-�F�|��u11s�Y�6N���B_�ⲇ������Kl&v��ˏO��F�/+0#����a�/��M��]�.6πgK1�`f�+������t��0f?�)��W���Ĝ��~+T���}k�ة��8�jB�`��2���9�N�Є<d��z�s��}�Q~+:u�5J�d���5�����-��r/�ۅJ1�\�[��0�*{>�_�M�������5�=|�i����~1���af�Br�(kX��̍��E��oѦO 8��Å���P�����Bm��(�������X�1�����������b�Ht��9�iE�\���:|�T6L-7R��_��^�,ry ��*��Y�����b���u�Щ4`n+���6j|�t5�ͦ>�6;���bz����������{m��Q&��H�z�7
8��bed������u��ԁ��l¥Kܥ^Tҷ�5�����(���	bB%�$�
�,j�3�z%v��Ln��:@���??�б��ڡ
�yP��)�ev{REG�T��a�]l`�`4�7�PzƋ�#��ԏ:�~h���df��w��~��S=	x��#�g�"ؘȖuH(#�c�P�q/�����@��3�	�c3� �q���gX|���%�6kZ�����Q��0������&	�����<dt�}t���y}�~ˆe�uy�Y�C�8]
�SΤ���_R���w8v�?!�(^�]Z5S�8V$�������[��q����!�@��Awjv9�(񕏦>R\r�P%��\�[8�mA��I*��У��K�A^_��+3�^����W���|쭟-��&x����z>��)�ŀ2�@���v!0 N����5�������C�[��J�Ou�:�o���H5���X8�Y2�'��]�L��~�{����j�Q�T)	�7����:�jXQe�K���YF�����m�+�kV�z~���tQ"2o��?�M5w��Z�.���~̞�{�H����ݎ^p�	�͇�>�$z߃���f�̓������<�@)s�/ vv�����B��8V]7������Vԯ<��D%�CA���%���X1�9�c(�՘����e�o��eLI�AnV �oʫ;4�G�.�?�Mn;�9�*�R��#�=何=<#�"�?>qpSȰ˫�j��(� &lr橡v#^�RW�]�����b�����Vح�Q��� 9d�A�����R���)6`m����Z��%kب��,
T	š��LT�(�KaCp�|�Ҵw�)t��;1�J:U�8�0<�S�R_��J�aD��o���q���:��U���)��#�4�Л#�E����E�x.��,%8u�S��7K��|�N�6fS��u\}�Ex��K�2h�ҳ��<܍%�=v�p���lli<W��u�p�
[h�"���+-a�;[%�������G�:�8
�~�n2R݋���T�Aq6�=���ȃ�?�I�|��믏�	�Y�:��%��!�fk����c�?�֐&�cf�-�5�-U%��1�d�iF�����fW�k��(�������\Y<���N(/g�[������'��W��; ����ּX����v��W��o%���<�yo��]g�V����R�Po��att��M;8 ��qEW��>h؆���r�����2m3w���C�zg9k�$U��.��6�R�f�`���~1c�E9ǌ��F��V��qKt�#j��iK�N&��Al�h��(��,��Bʝ'��^@��#�B�&&�o�?��W��jQ;D-]���8 ��N�iZԢ�w���Q�`�Fq�^Ծ����]<��3�S�����r
l�(����4f�i)��&+w���@��
2&5 m����)Rp�k+Lc|��(q�O���-B0�$����F��D�p��~^E	������x��|z��(�$db����r�F��AL�Zh������`E�v�`��.l�=*�ָ�ᐠcg�c�4��z�E4#/y�[��e��1�0cӲ}oH
�'g������N$a�p7Ζc.!�P0y��D:nѷ�SI�*j��-�G���n���|SbZ�iV�8a��P����9�CS��*rH]�~N'�>e��Nc���)�$� �`A��05��w��3�*+a�@�+̣e9�Tޓ����ͷ��8|Z�pc� ���6~�W�(�0����U碩Gg��[�875�G�c���d�8�d4��{�>���܀N�\z��a%dd�Z���~���U��$���M�_@�u�~9So]oS��7�xXS�9�8�+��~���&���zp�w����Q�TK�����Y"HN����jI=��0�e�$�P�5��U�⽙�d숾R3`'�.k��~ �����d�b�����隍-���)	{R1S��D�x��^�%&�vf3���QBN�mHD��f�HB�߲�f����b�~�1^ �abbG��@x��l��r8xAB'
k+�?{�jR��<4�R�]�zR�i������0r��F�r�ǡL�f2h.�c�A�e{HF���o�F�ϥ�=7�q�g`���H#X�hG~��0D0qC(�f_x���Cu�H����-��*D�w�D`�ٰ&���,$�@d)�7m�j�5�l�kE�4f?������Jx���{?��Sw�y{����G��s/:��2�FDA�
U�9O�}�ĩQed�~"60n���IB��cq�'o��i	SR�S���'C~������/��� '"��� O��}�CIP�Ƃg}������p�5�=ݝ:���ה��%$�H	H�=��>+�����鉌<�i���A'8�0xi��A*TT��H�g�gl��i٩������D����}�ȯ2�o��{A��+Z$0K��� <�N`����;�hӷ�K�i�Q%�)�X�v?�O�D����6�k�	�����#��w��js�
�����ӆ���a��;#=��8u�r�Ʀ��7���ɸ��5	�%�X)�	ײ��`Z��;q�RI@j�.Z����,�����y��t��}E�����|"�u(��39�>.�����&��0�X~�IX��:^����\E���E���_nnn�
rK��h��Y7�&�3f�c�����DLcV.��!�`�h6�>��h�4����?���\���v�����Y�.(hv��3	Y�0�)M,g��L�_�Z3��B��8��Uܷ<�3�+(�3^^��������:�}%�~#�n� �K|�a�gэ�@I:�T��vgSֳ���t�D����w=J���R�'X\1v��l����_�u�Ng��Cʮ�̏��}z��;(���o���7�vҶZ�� ��9���h�S�z���/p���	�gfʯvZ �f
��뻦&������=�ôQ�·��-킟y�	-N���'��}�1_����z�/��}�_�'�w0�Z��b86GGF������0��n�d���4�?��4k����k=�;XY���������8bm��0l":�ݭ���X�)�ל��-��22];�z7Fw3I�������PͬϨ
����B��G�Ui�ǩ��Y��	��F�%�K��0>�M�Z�`/�?ru���y�����Z�z����N?�f�.r��܅!J�-�5�{�Xx�[��,�G36"�|��	~~�/��6��_�xx?��W##��sarS�������$D�����2�-�]6k"P(#�f�m��[�����0�=0��{���$����R�t��&&�>���։�H ���bu���i{?ʫ�Ӥ����l�3:ZI9鵠;�z�C4����~���Qs��.�&���@��Q�l�H.�yHC��%��& D/���	��P�?���:9 ����\Y�+˜6}oɡ�j�hZ@5	���m����J�# �{��?��wJ��%2,��#(��"\.��?�>��!��]�Gт2�f
M4���%q�H£�1qˤv�U,�&d�oiP�B���Z�Y���㛀�� �����>���tY��Of��q���>55���b�� 0�P|Yh|>�@?��\�j#R�_�L�7k��W>�J�8޴R+�w����+�{xNi�xB�JaL/>|�Io5��H2vz)U����MO�P�/6�7?g�Z��� �p��p�j���)V!	Rd fFp��?����w�����2v9�mD��D`EgǚP�^|�`''�+�\�N�x�٤���~H��n�C�*���q|_sy����VFFO���v������ب%.�rFLө莽]P`z��+��M:�Ɋ�˱�P���٬������]m����6���YN,nU*X�x�ؽ��]+�(�C΀���/��~��̂�k�ݣ1���cvn��!�FQ�e���`P]��C����5A�䈓�OӦ��(���(֧VcJ�>�
��nm�esA�Q�͍rt�ŵ��	�{ew�ljW�s�<��E�G��O������EyF27���j�v�b����
���	�EL���z^_��0vG3�������~�)Dk�T*�i1FF|�K����`�01��3�Z-��4�$4�3��x���W,�l�� �V����a�g�'g;RhE�5V���뫒 y�&������*���J�g��W�y=*����X(��Oo��G���X{a!J�ƹ�F������-0�Pnl�]p�9G�r�qc���&Q�[�������p�/vHG��@ο:��zN;`s\�R$��`f&(������U��	G�|������A�����sk�dH�T�Yѳ��h����l�B'R��͖�im`2��`_\'��ʊ1��˭䀱�fŠY�>l�����ߔ���F�����(�˔1������S�#H��ͤ*T�Ȼ ����d�j~N�����S ZkX�!?'t� �[U14Lh�]413�������7z��B�X�;����X?7�����&��z��Bm.2�Wr�[�.ΒV���zz��>�@W*�G��w��g"6M�r�a�i� �e�����7e��L�Bn��D���ʩֱ|��P��:q%���щ�N1�T���q���E�)~9/��o5�pm�p�Ϟ@�%���"N�+��8�a_��^���~u���Ѻ�S.kE�x��経� �h��Q�[W���U��ce$���m#*}��ߗ����`�-��%�"m��[s=���!<�b�[�OY9�E�R�!� ,s��  bH܀��!2�1��g�������jx��a��5r�1D_5��S���j��ìL\\܍x���m������әx�7��>_����][54����gE�o�7I�5�ꉢ�Z� /k
�a=Ůڰ$?J�{�(]��&� Hz���t�Ő��*ä�KC?�'B�����(b�DjL��'��!"iS��Ϥ�'*��3�2��X�U�@�Pbc�%t�u�)�Kw#�`N���IM�ZX]���˫|y�8��9[Qx�Ho�<\���P�sڐ�1C���������f���Q��Kp��� =�/r�v�A��,�Sڑ�!w�������|Y3v�f[ږ
��rX�\�h-�S8ևs�rD:9 ;����([]����hl3��̡�����nM�p�x�zo�v>����j#�R�W]�)m9��Db��	�sN��蕚��Q<�0.&6�GN�Ȳ�Ϥ�����Y*�
fh��DkcK�y	GG6�]�999�2�1X����G�~��L��+��Zt�������щ ���I.GGG� �f�7bC�t���*D�xޤ��L���/*���dѴ���<=���BCa"8|�ӂJ��YHt����5��x���O�e>w����lcp����)b�Fp�DKf�~D|db�4P�쓍�?7��4A���P�B&�~�#a�^�q�,@��䢊�f8 \`nn���ڽ��@ӎ�U;Y�E��6׫�b���h��%�hj��Gg0��__�X9-�Z�����kT8=_����I<�j��n[�a�����>E����lQ2��h���lV��H�=���Ÿ�]	\F�p0���G��=\;�Tت^T Y����r���ݯ���&�1@�K�����}���#��]�6��&|3�]4��2q�l�k`�FE���s�yH�&\��,��:�hli�l���m��!�-���ڮa��-!��Hw�� ��t#���ҍ�]��i��Mw~��z��C��Pֹ��sE���5�F�33��R�^�&�!�ٜ���o]��*B����I���V�B�u)��d^A%z���f���Jk�D��ν�SY��B�Td�r k��쎑Q�bx*��2��`��Z��v��8��_��BY�Թ���Z�p�2_K�=���{����G���d�o+��\����a*HK��zg˾VYLѴ�nD��3�
���'��=9����oo�oDJ��y�ϳ��}Lҳ���s�YAMB��[W���4l��ݶ�(�0?����W��%f�W �"''��X�����`<4d�勥ا�Թ@��Wʋ�s�����	ּmq��Q���*�G���ŶE9�[�{0�V���_�E!�y�YD�R�A���*�J;��m��rm^)5���H��ތXd*���]}Z�ԑ�9�/}ߗ��a==33���p��Mt6�Xaަ��6��?3�U6� ����$�-Sհ�*��KE����'撴�#N!Kb�gL��j����M���0�đ�m�ȋ��Ig���#W�@��nP�'��A��q�ۙSd�;݀Á5y�X��R�f����~���|I����=��$C���_9qJ����hMԼ���d�Ywi���84$�x��'6��I~{��"M���)��d3RR�ْF���%�����Ȗr���@���a�g�?�LP^|�%����K2�����K*#ww���Q���xm���U��p��p$;��Sp�z?|c�K�|_�^�d}}Q�Y��F��2���nw���R�Pa���a�/�K"ڽ'�]�5[_����>���uCT%[F�F�ݿ���f���3�i�|���F�����&?ur(HduY���2-��X&���(,����'�C'���Hl���O��W��I�-���(E=<��AUm\BWxF+,5\��b�
�[��)�FL����uk�͇�����9Q�2������5�s5��5�:5&��'�ĒVlT9��l�/p6\0��ب�Ă���(j-�1�-��c`��Ы��y�V��;&O`���[Q�r6��M�NQh�������*���@]����j�)�J�J\�����fx�_-(�Ωm���:p��[��Nn֮��e�^ł��;�}E���]�ll5�pr�`Mm�Q�Ɲ4K����vO�Q��a��=����Op��}tq�\��%R�?4-�2��f�7�*�����b[!zhhG%�7\�8�62ߓ���L����q��:OA�����ֱ֮2�v��훹�P��(��r`�}	5�7���<I��BC�l���9�Ρ
�e��zS�E{H�\^K�Ͳ+٣��!3��aһ{Y �s��QQW���mK���9*֨���)Tb��0�{���!NsɆG�T�?��Y���$êx�-N�
��À�NHKcH�j+VN?R=�o���B�Z���ұ�鸿�\~6{#vP�o��4B�#~�+ڽ�/�ʔ�T�?-��*#����{��?b/����+%����Mvӌc`Sly�Dh���xr~>��p�gY4VvX�l������A����D��"�O����������s����
CKY�|":4�N)k5���aq�ט�v�0�R���i�_�p��z{(����°������T*��h�C���:�ۿ-Ҹ�9�x]�ǂ�1�,��_�w�{�:(�Jٯ���W1�TC��AE�܉��l��!VA���0��yo�����SR<k�����P}��d�o/!��u�H +=��r�5�Hݤj���V�|c�j��dD=Z��{��^�����K��G���S�~f馾,#LG��G�|CCJZ�1�"]�G����h=�W�����(����?�����Wl�����Y��q��8����%���$4u&��eml�>��^z��G��|��$W},���:}���ձ�9�zODA���>R��'��x��&�a�� y�0���-��}W�+�p��x��Y
�Yq�ڙ�	k��8�2{s�'�T�P;/�����ϖ<����7bF���5�Ι�fPU�wQ�g-��0���1$�u�gR(�-v���F���{sYD��U��6�hʓ�Uu9!��6lE�䲚 7�H�O�2�����[x�k�jDP����'f�������r�
�mw`�y5C�:�9�R��'K����L���
c=�\��R�O��n��N���^�&z�����7J�t�Г`�A�"�dq)|�o�Y�\M��Yt	XM�A����1ٜi��Q'otDvw�P��ʈ_Ζu#�y�.l�A���?t��!-�	d����"����KP*����w)�㜬��0�����``@�Z���5��_҅���S��Ư��ğ�\LX��H����+HR�b��
	�yA=V�XAH��pz���'������h���2�C �������L[���$*�Ac��B�Tє��J����ug4�l�(v}���y�D����1�T{����{�)��W+�����(����v�o�9j�ϖ;�����ch�`T\���.����Q�y��e~$'eP�Z���瞺�����w�bY�Q:S���
\�v%�T�sRW��g�^��GO�
 �3��Ⱦ�/��^��{dU4�#���g�z�ՈL|"qB[�7�^u�'17x�ј�dC�(]���c�cX���Th�R^���nF�v�rN)��6�q�����͝���Y�$|ߒ*o�`L����>���
X�~����j�5�	u��i�N���HY]p8�I9��?.��®�AA����k��H�P1��
��Ȁ���m˛����o��!�����h��)��tI�Ĳ"��E�6x����W��0�����G��EF����Ʌ�����s��%RQ�)!vW�&���:��-R��I�K*\�)��b�leM���sz�B�f(��,/�ײ� &�z���]��b����n؁/�l����մ|0��ڴϚ;�j�C��:����:���|�
#5�nh�������gZ�E��bU��$,��%�q4�+��F�/^�Ew ��|�B��4���uW��(�ę�ۧ��u���F�3dK|���oc7�/[$]�w���Fg�w!�v(D/�'�o�嵇��(۪+	[��$-CD�W��4]X>Y�h"v*♓;|uV�<�%��-�,�W�iJvv�5�)*��V��7�Q��'"� e) ӱn���tt���t(��ө� rc�Yϥ�����1�D7�ĉz k��v0�w{89�d������2����	+�$%�co��w1��WW,|=�����#�a�kL	
�Z�͉��@�._"xd{e�y��G߾)2�|��􇨼��Ak�c�gA~Hg0�nXs3?PjGBBB��%ةz������p�f�K������a������E>�z���\���Ѥ3�������G�)���3{nͥk��Hz{��TipDD���èV�o�l�x�`�&�M:�e�F6�u����)��Ed7��0����\#9E�X̔L�Gm�)Z]�N��3n=<*���m�1^|�U>�I��f�G�0��V�����~�}gTI6ߩ���}��ۚ��\61��<�=|=�H�0r�I��p5�2�6#FD�k���R�'͍ĵ��ROBBH������g��P��T��{?������%�GW��G�@�%/����8~�'�'ˣ0^��C����~����D���*��I��1q2��(ގ`�:��r���|i�LD��쫃���n͉V=GA>ը]~T�p�͖�dȸ47�E���� ��2�2�!8����!q������Kt�J�Ԁ�mKo�Y�*��|�O+E�`9W��yҊ@o����\䊍	���?2TeO�ДU��b��I�<���Qu�r�`
�]w��i�$��g���F|���ϔ��>E���WF���	��~�DQΤWXlPN�5
Y�A`�N�������Sa�� d��!��kj|�=n��ӻ1�|>l*�t;��H�9�1�pg#�4�r��'���ZHb�ecTmЭ�-�����M�,Z��ap\E���>�$K�~+Y��ѫ��'>(�񉶥�������I��r��L�.���$m��+��{��cΠ��ǝ6�J�����}��F�������v�N#�wz��/*%"���Y��1XIOOҬK�X��`�C�ݧ2�i4���:!���[n����h�	�؃ϒW�N��r�M�B�0ޣ�]%չ��p�`�|����8q<c�/[�P�_��ưP��~��7�u�A�#���q߃&ei�^�%?�@i��FN���������F8-�!uXS��<o_�#�>�]�cQ�E�r��������aHL�~���>_�
<������ W/��pԨ�h˴y� i�lon������꾫�Vv%�IҸR9i>�bF��G,�eפ����XE�S�������MJM[��6��%�����ֵ�X���>&sO���������3wJ������Z
����K����O��0�/TG��	Жؕ�R�D!�1+?M� M�QP}-�����,{���;<�f6�1�|Ԣ�2��C5���s���ۓ��÷�K�Bi�(*wͼ>2�_�����&8p�ս���ۨ��r��~�) svv�Ȫv뱔S㨫��΅6~�=l1�C��2��cͩ��`�vr����4��I[�Nx%���=@m�df�T�nhP��u�]��g�@z9ɵC�Rbe\��w�>�ٶ�?C)�m>X:H<�o�5c��ÌW�����ۂ��c�7���F����Gd	{�:� ��qy`x\�Ƈ�����yf�l��}s�x�{�lڥ}�}�}su�Q��KE��;�����+��������Du���f4�B�ѣ)��_M:ϩSK�2��F6s����p�dd۠Ў!��v���o�7~�H@��Gr�^�O/k��W�%L�~s��ߞ���WE�;��}_��ƴ �[W����+0�:K%4B�X6^�f�{�����#Ô	6nV%�W|}@�o�;Ψe��/#/�a���l�VE5����\���j�i��3OG�;���\6��S���j.2��u�_�/�����w��@�i�n�*Wc;��S�B��[E�X�����vwBlvw)��#&�Q�%��l���{��3{~��;�vE��۟УRNm��l��t���τ�~6,�~]c�{yA�5���؝�3���}3�՝���>����d��|�G�-
�! ��']sܪ�&��@!Ш*+��V�8����e��7vk�A�+$��F��&�H��<�mݠ�hE�W'��P	�n��ݻ˔�}UX�"�t����8�E�-���B5�M����O���g�@O_N�(P6��C�CyʥDX�y�^���
���v��!"u ����9��MOOM߷7�/7?P��G27f�F �p��Up@�sj��b���FB�h��.kEhܹ���dx;�t7<�4�����w6˞��Q��{.��Ĉ19����|\�:��E&��DL����>�=�S�p9�X3�+���8�1�ڍ���<ߞ�	~C��+D��֗�pz�$���x����ߎz�[��ټ�A:k�� pg{#��(o��6�E�CPUd��,�i`�u
zS*W��4v��_���˂���MT�&gf�ّ��X�9�3j�d�>�ܝ��l����%��	�Gy���x�6xG���혁O�q�u�ȫ[84�	�rrJ:q��Q��x@f��d�����	�$Wn����%ڎ)����S�^'�n��L��-+���:�)3�idE�!)˺n}Xn�4cM��4��di���)�	����.��� �-�ק��lv���^)�ڰ�_��$ �/�)]ۚ���VP ՐׅT�}���n0~ty5?�a�F�vye)��A&�o����N0Eq?�omoǡ| q�M��jXv!�fi�Aɟ��/��z7��&�~p����V5L���-�Fa}	�o���bɋ��18��S'�P�������k�׬��d`��*��I,�u$��<έ�]����e+��J���7�3k��J<��%r��X���p����$�e�⽢Z�6!ɉn9쬶��4]P�b�������7�h\V��q|��·=�D������x��y�ײ���;J@%�С�᭠�,ٸ���ڄN�c����9���țm�/��������N�i&w�i���`���gՖ�y��@��ƛ��á��?8��(�o5V�\5ҩI;%#㳇!��3���GF���}L<�a�q�G!��pE�'������,�D�%�I�z3Zw�hE���X�c#������0���l���#�D�:��BK3L|��!�DR��*|i*����71|��� i�VZ?�'S�Ղ�/V���� t��Y��E�ƚ��#���j$��$�V��2G��~�(g�����-�hU���Ig��������إ�C���_�)6G������o���+�-��p0��xYUx	�x�����XZk�U4@i�ڙvd�6z1�4Q�Y�����#ƐI�~���)9����o!ʭ���.)K�#4��%�_��
�w�H�/�P�,��@n�*���9������,�q������4\ ���S�©����k<x9+IˀґC���3jk���� ����pr�7��g��y�a���ݥ�o�g0�q Gd���u[Kl��*��8�,�q蔑�Q�T��ˍ\"��I;$�H���s���-A����@Ә�!��j�&��5`E���E�D�����_�)%ipp�F�!"0}"E|�3. �V����rp~_3p�C��TE%26e;[��7K����y�ڛw7IocW������C ��~v��J#V���_�W������YBV6~r�k������+����(�&K$#��-R��jNY[�pb)�r(� *�e���C^�zݲB��.�O��-T�::$ ��:������>�3�eYx�6xW��eV�������^�M:��MD��1Mp��e�7�;o/�@S�na74v%D��9����D��x*�P�L�S���l���S�~u3^M�1��Q���Կ)Q���v������sO��-��w��
�t�U[}�5�������:�kX�z#���s�{�&yj$����4b��b��ܴz�%��4�K�B�@�-Eķ���Zr�@KQ���҆��RD����N� U�y�e����z��]������}q�K=�DZ.?/9�VV�z��X&�~9�vۋ����@���0����-��^ �D��P������ɷ@O::Y��~b� �Έ<���oH�\M��HYk�� E�>w�z�"w�·k���LG.�LDL�Z>飦Me����,��|�~�!�5�a��2�- ^�o�ݿ)������������L�t�p-]�m�v��!�Bs*~x���O�PQl��CG�J(Mm�&�\��\�[���`}īt{C��	�;&�0R|�bWO����c0�htwk�PZ�T�\��P�P4��L���ח{q��'��z�њD�{��9hEXI���d��a�ex;��WM�5�`�̖�6�t�_so�j�[����H`T����ͺX�F����k)w�e>����tpѤ΄�(O�����+��]��ȴS�s$v��{�^�q+��uw�x�F�M:2R�"���S���k9x���Ǡ�z�c���%���5E�s�M����}D�n34������`$^U�4��1�(�P_��k�M/��b���!-���w'Xˢ���1�3Y�aĨf�<�p�d���c2Ǝ���"�e�`F�eI�i;��~��h7s$~��ar����e	2��I �55��v�^ <:5�:K�갔-��'AC��--r��D���
 51$� � �{�F˝��ů���s�z���t)Vn]\�����}fk��o��/pm3��VV�i܊��t;3\r��JP�W��u�dϧ���@C�԰�5r9�QNi��Z}r�k�r2��9����[���i�ZH���Ϻ�9~�n�c���c3	azϓ��B�-3og�������+�j�����>�}��g3�(�n�KoC=���ݴ�kn�a�z���V��%�w���5��|;�&����僋�$c��z�!��e�TOc�����7���G.�_Omu~���mm���B����"\�����T����-�WF`5ޤ��Q�=.���D2�~C{c�.�;���:��b�PJ�iE�g�C.�.��;�J�K<�|A��Sf|�To ��!9
r���S�A/��tI<&s�V���&���ӱ��B6]���="�g�J��<�@�iL6�iy`��M��
~m�"<,�V��f��Ygm ������M�����z`&g:
��$�����?�C����rc��ܓl���y��y�V�4�C��x^��m�|��h��1�sR���*!Uo��I5�kj" ����W_zy�	�
���v7�b�>�=�/�Du���+����T���ۿ���Ҭ��)���]����,���i�[)�_dQ�+� Z�T��ifό���ܖ�XE�����T��k,�c�ǿ�������?,k���F��C��_�5 K*���4�ˌ�RG�3.b�H2�S& X������o��
G���`a�*����0@��x˿���!�����������-�2���?�M�7S,Ny���#��춏�R��r<O���ߕ䬚���p���n�g�PR�j?"�d��v�z����HcŽ�QAR�[<�}x[�|��: Q��ܻ��x[9�Y
p%e��(�%�l�8.�G�9�0b���MQ�N�r�o�>{��D�JmLczY1��'�> ��+�7:�>��4�v˰�B���x��N7X:�I(�q���`�K�\0֏�I'�绺bخ�#���?���%n+vǏ4a�.��fS��U���?�mT�iE�$a�8�47�������N����F��;����ᴯL����Y2���߸#`��
�w_p�>>�?+���x1!��������u�l�n�3!�"46#�x*jWFW�~����X�Ku��k�1��qͿ�k��LhQ��nN6ޡ����z����a��k����P�Yo�$�I�ysZ8>8	;��o���e�ܤ�ږs�)�s�W)M�`3n��^!��	�Zi��sc���3�av}�r�k*��+H�wk[,�b[?x�6��p6�*��
E/4�����:D#�A�K������q��[-��P�n�����"P��G�����,��(Dͫ��Ȟ�i_��R�W�i֦�2���E�XD}Ʋ~��D�F6�\h���2�n<f�ޞ�9MSɪ[idj�yE�+1�N����!I��>�x��G�e��*�;���k����gQii�(�j4~�|��Ag_Q�?[.fs���a��ĳ&28�U�f�ኛOK�5?��Io�vv��R�E��o^�h)��/��d�{�k冚>�U�����63@#�1�}>J�4�/?�WS���ͮ]+�/��\���x{t�S�s�$�yB��s��"ݯau�s@��l�W6NN��n��m�⾛_�«r1H*QLp0��ba��;�z�?-�o���ƯO�f���-���?���ډ�5�hoy�9%����V{w�#"O۫�q��A*2($�c�1I�rWv�w�x�������{3V$��k�H_���_�T��?z��=ݘ�I�@2
��;�����>���&�LSSfo��i���Jo1j�#����P��S�Y�w*�����|x�'�h�+�/�+�R��~�[f_�;-��-Ҏ���������ƕ2I]��~~#m�i��v�nk%�د�m�����e����g ���fY��d�Ļپ>2����r��5K�����[.������~�%	#
)zZ�fZ{5�b�T^��V֖b��pH ���oȼ��D�X�oF�T��jxЉ!p2�^��k9ra3E���^�4Y�~2��`��{p���إ%mm�e���?��	�f������#h��f��g�~d5�Ȗ�LϏ�r՗L�����)2�N�)��񜭞�E`aD����m~�c�;�z�?�v��jf�ǝԩP�G��cW}��JƬs���dt��7*�7��`���w�J\���x�)���~N��ӓ�����M箉������˩E���GZ�>FFT �6Z�ݮ��_y�GGz�2I��f���!��� %w�b�Q�P��7pU����d��&Q�&n���`2��O@f��p�e����DC��D�5���OD�g�1�����+��SV�GG��.����8�A,��	�ۋ��[��zӫ#�:NF�RQGGGe8����:n������}�ߜ��?����e�����H���mhÜ@�[�N�_�n%�ޝ?X��NtS��D*�ȸ��o T\����� �o�Ji;�R'VUS3u��l��Wb?
b�OJ3��&~���z�L%���/f'-�0�_F��!_^7n��!�t����R.?�/�$y�fȹ=�~]�.M��U�G�SD!�أ��M;v%?��*��J �Q�QS� ��5\d��H$��]�}�:�%�?�y��-�<@x��s���c�؁��B��3j͏m���\���Z	ږʟ���l⵬k��H|�L�%�c��x�5A��}h�������ʉ:]�J��s
z�p�D~<ͺ��e��M[��:��BEaC_��Q@���P)�&���w��y���%��1��DKS��,E(��h�&���_X�{:�-y�!A����tkcD��b*��"plL~��c��Z�7�.+0���.���Bb<�Wyu��7�A�qAI?���_?���|�c$H�h�x�]��~���l�xX�Q�����B��~��Y�,� V��6�#͏^Sc��%���/�ZC���J˅��j���=��TE�(ޑ"-��z*H��,b�����y���Mz�����e�b6.H�ңdcL�^HKj²F�L�5��ƃ�]/��[M���o�O⪿7�K��9���f�X|������t)Ywi�^"}S��,��"d�uq���t��a!�Ґ�b�\i��&�M�?i��B�ܼ�m	z�Y��ۼe����!�:4�ϴ���^�d+wji�Hf����.���x:�.�tE|���-9����l^������{�v����� �����?5H~~z�^�+���?��k/��`��y��vC<�s������C�6KWVQi�1������G���J�&��h�L:ބK����-�-��I�zL�w2=��D7�/��� mtnW3��P�P3�	���7hhhvw����:ff� Uv�LP��"�25bb�q*jQˀ��V�jОF�k=���4w��~a�~���;$��+�W�aN�\�)��Ĝ|~�&�m��7Vz=���I���K;v�W�o��
7qi��Ŀ�{�͙qE��>/D���af�j�l��Z.��_����T^Pm��37`�P{C��}�������FI%T�L�m�����l�䵶v���Ա��Bc�hĎ�~`����*��@L����6�QQ��!��3H��\���5��S�P�԰l�spx��v�� ��Ll�X"���p�Im�&��������8e�	7t����v�ł�e�:�"��@������́� ���P�.��!�*�q�`yc/�Γߩ� z��A���K�B��t]��7/O���n��O��2�)�%uL��V���.R:���F"ΐ̿���|'KqS9C_�H��6Oϑz����C�J�㢉���:�o�[=������\N����a���n��k�%ԊB�r��ףݐ���o�f�v`]�$�u��Y��$�F���I� �#��H���XG��<�)5��y�@�v?�mҹ��D
�N����3���B�*�����dϧ�-�-�1ҧ3�z��9~VV��mQTU5.��q�R3Z�ˢ��UK�Q9qqT���Γ�y��V�>�k�-3k�[��1�;��n��f�g=/p��[�^m��TM
��,YO�����0k-�uE{�Q'+���@F1���ɬ]�'s�����Q(�F��`�^},���f,�V�Y�z���&ƳŌRm3�Ums��Q��,;�bn����m+N
X�f8O���8ӌ�ͳ�!Ɗ�/�:�W�ג�w��<��P�jߖ+\ﵟX��U�l%�J��n �������7���G�[��~T�\(�&�N>�u��\��S��^�Iq�£4�_#6Ȉk�W� �=ڌ��ǒ��ya�h��>��B9"��J�PL��<�	 ��2[o���^M���GCn�ċ_5
	�ksRg~U-K��_\�W	�dȶX $�y\�&h����N���Y ��n�v;o�%ux\[G ��I�瓤��N,Z�m�� A��|{_��jC��ZG�^T
���D��e.�`q%��
���h'Tk�_�"?�0�rդ�=Bd��9�m�1|}�'9jU*d����8@.��qW����?�B�kGN���u1���Px�?ؔ��0YI�{)koan^`���o�e�3ۡwW��-�~��߀� ��AG&����V`��I�.8If@��I��<���s(�◣��X��]��a�����7���P�w?~�XK�j��t�����Ω�n��93W��6ǾQ�.�۵W	���.��-V�K�-9�00����"��s��x�C���]2>�[��ͼ��)I����Q#��-A�^]������
��J�Y��ۼ�Y1�٠x_��X�,BrUDU���!�p���k���i%�H$,��=��,n'	1+�������PQCp��I]]���W3@� a��>���0n�D��ʉ,1���-��qCj�wu�^X��5�^����,��~C.��7��ú�o�A`9�g����1�}�F�%���ˏ�tZv{�$�TUy��g��?Е��7�	��E���gy�v��'�տ7��_q�AI�G11��>�͙c5�4�5������)�u��l,�"�D������b�{	�]v����Y�;�y&��{d����^�	��{��j6��*��.'9kxɊ��
8Zơ��h�`S{�m{�;
�E;��Xx�4�F���>G�Ӣh��{?p������n�^�G׾�W̯�/���p�ll��Y��'�:� ���gT���,��e+iW����f�w43��|b8�^'��N|��9!X(����Ծ[��Ӎ��܏T�yC��Z}�`���R�Gw��x�q&'YD*9�d�̥����opc�{�����ٝA��ʭs�.z��Y�r�<U�\�럇�xxF��g��n���k���o'�L�b���`��y�Z#�P���E;R��Z����aP�c�W�B��Ph}�m��>�ڝ{�!��Ɔ����6������	�޽�򪫕onli|w�⏫~g�1�3,�#FW�L�{r��tnuAr�lXʏ�M���u#���3F��~f����f��`���7��K���;�ߚ]���C����O+�z������� �8u�xc���Uc��R	�l���hW]���l��;��j_�I;<��a���I�`ʠ-�y����pں�%�q��ļ}��{�g�:;����9熪�Կ|1�A�&8_k�@�Bh\��P�V�:��{Mۯt2�iU��v�w���,��(��\Ri+��~v	�SG4�J��-`R��	�����]ն旝r��;Ocj�2W�ObG�z�Z�lh��.ɯ�P@2���׿学ԧ$M�����ۺ#s����C�F��I���NZ��6(h���6x���s�i]X��~�2Z�`U�+�,0y��5��m�l�|<�6���"N)U��H�?4����șc��u�������R�l���]�ź��ރ��б|���7��:vk��m��0�T�Q��y���&C���� (:���-K�j%�PW(�v���ۣ�jܝ�o�;�.�>	��L(�4z�x�[#�J&4�G�����ɜ��}���Pu���\��M�.�����e\K��
�Kxy��8�Ɉ]�!��q��RB�#��x�]�������s]A��'m@��`�� ����p���̿�ڭ}������(�(gk^PSg��7]~������5^e��h�(�.���JY�ݹY�zo��	q���y�s��-D� 2�R4�!K܄jz�|B�W����W>222vP"��r1ֽ�}u8��Y��Aj�������% 7�51���*毴�׶�U*�+�-_#B�eׯ#l4V4�4�_Q�s?ּ����j��g��s-����Y��=�p n�3� ��Y�I�Vz�%�Z�������^���|#A<ߩ)l�>�s��g)j�P�ܰ�����&��4?��?�r�/#S��>[�����
���5I�Z���t��������;�<r��w��#@yꎳ��w�I�K�}�T��k��>w�m7��'}�:� ���hXhYk1�כ-st�V�ش�K�XJ��ҭH��S�u��E�ZL-ϐ�=�5E�q�$�#��Kc�["|�Y�p��F+u���)���)�q]��w�x�̧J,��,>s[q�*�z�m����yI�j���r���s4詄��p�� 6*iߋ��V\R.�����0aj�	䥠�#S�Ma�(Ĥ�'���0u�h�i�i����u`1�5�ԍ9�s�.���v�C�t��v���g��t}Dd]?�T�w��]��{��@u����ZJ��}ȶ�<�Y/S��0���@[�!2�˧�7�<=��"���1�P,�%f�rHL�.���'囗�>���q��u�O$RPV��c�T����t/eQ��"�Ъ�Ҕ��ɂ�_	ǩz��1+w��,(R��L�G��,�Q��7�2���)�Mv��� ��!�'����w��O�Џ#�b�(t�r_<~��s���3Z�j���z�M�8�ֲ����.?
>�nSԫ�ok�ds	I�{���s�8���WM}���q�L�r��*�G�ƀ�"N�w����WN�M�F�JP5V��V�̃s�v�^^$�aʒ�˓�p��@�0�QL/�,�������ː�h"�[Zm��hN�ۭ7
w�{���i���թ��	�O�!�_2Վ�y����B^Z����[LٯI���W�(�]?J�ɕ�^g�v�EG�v��i>sC��[�R�Wr0Vs�ʞQD�*a�0�ı.f�a�UB����\�A(B�m�вݠ��b��|h��q��s	]QJ��HΩ�e�t���t!<�����f���`CO!��,9���oH��>�-;�[��
�eEٚ��3��5�ب��Tux��k����?`"�ݨe�.����Mb1�L#j"B��7�+?�����q2���My�w� 0����/<�4;u��>;�d�a߬x���Q>���걞fY���������J�)#ݣ�A�x�'��0�a�t�V���G����'n�����w�x�q
�ە��d#O������ߝ�m��<�"�8/�_�@��u�x��],D�����coF�=�����Le�"+^�?oD���m}C�z�W�1�K���!�@Ϻ+6l+����P(���I`?���K�ͬ��u���,q����1o��]��' ����@��3��%�U~!��B����\{`0
BW8��[o8���QmQww����a|�;PfZ�W��8�@A1������h $<���DC��<+2}���kh�N�<5����4
��d�P���H�T�]�Zq����C k�J�� ����f9��z���w�JU�t��-�~ �ӕ		�z�5(&�K�[����BP޴C�#9�L2�z�xx��BQ�{�Hg�X��� ޢ��8O��7V�d/����:���Q`g�`^�����=��A#�T��0���mՃ�!]�'b'}���U]�fީIO�s���Q�KRc����s2�U�Aʯ��}�'"��<���"#���z_o��WEb��C3�pť��M���J,)��P��XK;��Sl3f�6�J�PH+p�<�cp����{�Y�7$�u4@=ojյ��h�҂�N9!�k����ݡqzӕ�T�]�-��3��튲�T�3-j�����a�,�K�������t������KG6���X�� k���p�b6ƀ�sR�ˬ���z�V]��K��6#��ф���x�M�Y�����
�3m������Y��=�TH]���y�څ�d�2=�4�ғ��6�fD�~hWⓉ+�%�(k'�4^m�%M��D6�\a���0��	d�N�J��k͑$g�X5
�ݞ=���-�T>t��ǩ�����4��_-@�ɇ��
�Ƌ<��6� �n����G��G�B�PP���W�ܞw[�S<����q<+<5FX�H�����E|w���9��ef��!>������-Zޗǋ��n���GZ�5_�� �Ʀy��:�!�����C>�X^	�;Zx�%u	pB@��D�yi6�X.ő� 1�s�Pr~������0�?�v��-�p�c?��=����^4"#�`�0�<ã+�:����k��_���])�qb�5�O�䕆��0����hj�{iT
�{�n�1�o�;��G~�`���C���p�~����P-v|��jQ�҃�DM���@�=�1F�~�q����fw�Zw�i�[z��5)]�7��y��3N��)��E���#ꭣ����q@:�� "�ҍ�tJ��tץ�A�����N�KHww�����~�\ֺ뜽��<�̳g>��!zz8.RZFw
ؚ���=l�S�=~�ؤ���ViU�o�(��[����Z�g���65���ھ�?c����֨i�$;���K�����WDxڷ�]`�<W!i��[��o�o��9S�q;�P�0)�Wz�#��j�#���YA��$a��0b���M�{E"6���&K��Y��t/��1W�tɗ�FbU%�����)�C�,u`���
=>������o�)F��cKz�ڰ�ȶ��d�	�g \��� _�]�n��X:��J�����_�)+tc����S�ɪ����Ah�x���dg���]`��R�1�� �B�G�F�������T��0�w/U��g�|p���,
��b������`� 益��\��7S5TK��QȂ$�>����D�Z�ϻ�Q�a	>�ɳ���E�i�}��'����%fWa��,{����`w�(kDv���	�K7�Ph���޽���A�^�%��,3���6UA��Q����^p��ڞ����L�iJ�j���Ep�@~�A�%q�~�Ulls�7��u��t�T�(^���@x�Ӏ�3�:�nz��`�o�@���٩�����P�(�NM��3�\���L UpvfE�A�i�5����sVK�@��e����0��;�I���g���=We9�U ���8S�Y	��X�/5�'�V_q�p�v�L�|Z5:��s�¾;0��8x��~K�����y���Y�����]���V������?u�\����@���������6Q��w>R��\�x��\O��J�iڻz��k[���0����E��?E����W7�T�2K�F��cN"Y�C�%�\2�Y/�^����Q��UH��1s��i�?�~-z��E�{���w��*`�l�W�_����.7Kl��B��J=Ijj����|���Ǝ�ǖ�������ɘJ��@�U���N�p���d�ˉu
z-F)d�v�{��c���F?U"5�c�wZ��1~^nL��#B����(�V�T��:bOp�fdg�-�[� �0>Y��ip�l�������
���$���}P~M���*��d>��C� ��K9Vi$��\kS��6c��q�A{���&��ǜ��<�e6�މ�ы.�ĥwgV�t銲��GaFҭ��=$�i-	�+�+1��p��R�>ެ�oɟ:�8מ���F����l~t��?�}7I�����kv��p����x�4��a�|�c���{FOI��h�����%,��S�gKGr|�x�m�me���W����h��?=+��j�t�&�{f�}��B���0Qz���'*�EuI8i�f
C����0���%���j���L�>lĈ+��@�xS�'�
&|;���5Cy�9�+:>.�2z���w�=Na	�K��;PDv�9��_�E��z'������E�O!����.y)�`��B�~� R����E��ܠ���D�\�3�e��}a
l}�$��C��f �]�R����=�����ԯF0cv3R	�_&7u�]���Ven��Wp�찒�<�W��:stKR՜���C}Z��$��Wz����v?��E���_��?u�}�|9Ϛ�!��O�׶��Mnz=E�;u6���ֱ�;컨ٳB )3�S1���|�Z��ˣc8K�2i�e�k�o�&�'����ir��oS�}�lF���`�ɀ�a�2w�`�}�VR������jة�w�W�m.��a�>�o�R �;;>!�d��+Y�_$""�����F��_�P�x���P�L�-���kQQQ�k����c6²b���jf� �V�/��ퟛ}8z�j;OF��b�7�cX����������%�1���;���ВXO�A�1�mZ�������׼�1b�6�}�M�|��9��6�I��0`�>��W�BYNm�p���HE��l����i댒�Q�O��*"i�Ob��|��k�����������Pii��ь�
l��e|f��	�J�Ji
7"���|��(~(����UC����܈��������E�����e`��
��^Pцr��	�{�q| mp���m)����a>�U�t�~ӱ)�
|7VPLd���K�E�������CV�(.$w���>�U�@s��H)e���$�a*;$���N�	�%��^
�rh)Ƒ�g(�����@�����z��i?��ؘqѡ���1����֙3F_+�n�lti���]�=DCMm��I< v0}�R)�\{|���?5�4�C�qؒ.���'S<��ܘJ�N�]���cE���2F�]�s<���^W��H
FTL�\k�	���,�|��+��$� K���mi1B�ii~>�Pr�뺂�$pf��G6���A�iȬ�FJ
�T+��`�n��vzMU&")���/�\���L��#�Jd���o���<�ҷ;�!y�<D"ya�'��T�qC�&����C�bF3�����&+����S�G���~�!�/�h�H�,�$����Z��|�kz_����iX;��b��&�ƪ'E�=��x�4��eV	U.��mQ��̗�u3��K����=9m��ߔ1�Z�p
�4(��f�Y[s��`�X�h��-/\�Ea�jq�� ���4�]`�S�k�M�?f�Y#Ѵ���i<g=��%1z��|,>Vk��X�P�>�@��hAj� ���b�G�U�������ƒ�9��ׯW��.��γ�w�������Ҫ��hR���P�\BBB�����o��&&Vu����`X H���z[�]���^���}5j^��8����|��U����M�ý���8&���5�Cw�Y�8#F?7I�7.�1DXIQښn��Gy�4�]���~ge�S둌����(��"����U?��b�����9�4��&j!��nu�[V}4	�$J���_H�H́���es��8�l��<�17	TI���[[[�}PN�䢟A,�MU �K��$>��D�׳���)@��~��d��R��VY��*S��͠��2ER��Ҽ����9��\�D�u��n�̎�?A5�k+%+�/G_���K���a�/�L�c���⠳R���GU�;�ýB9I� HUW�����<'� @F�����*�������Px¥�ځ:�՗wW�<3�A'k�o3���c�̜���ol.pjFC�oC?GT�.��L��z���^�=86\�a�W�{uE&"n�X#�8��9�H߄q�5�=F��ڳ�~���]�a]�E���z����)$	��X���7P�����g6Rw(�x�\,�av���xR]�� �o��
D� ����+@�*�H�3�_��kp�˜x]�G��RӬQ��s�p�hr�{UC����AU��~��d�wKk�����m�K2��s;�o�>��|�#��6|�nUg�iv���@�'C�<���Gg���d��j�n���]M*��iϼ�apĮ��f��}�t�
Q�ZA%��b#������}��0��׹�kc��>�V]x����*�������ժ�m�ݖ^S[�K����丫� ڲ!k+8=|��*�Ę�:�9��3����H1e��$C��8�8�q��f����?��*F��پ/������ջ~��]C�����c��S}���2\Ҡ"�bSF3�5���DE���>�-��	;n4�ݭa�eV��^�n��5�V%D�9��� r�|�M��Zfw�Y�N��']�:)�+���y�Ar1���;I���E���9+ƛ��(�z�
����!a��e����n���=u���cg���jwd�ò�_�n7YЃms�{PG��G�qs��Gr�ˎW�<�ʏ�����£*�_r��Լ�ڻ���2 ��Q��Cp���!�&$H�g*���
9jW!���Լ�b��+Y�
zuU.F Lk:�<4���&����e�6��g�	�}^O�j��`*)Cc��.YQo�����2����}�OoKqh)�����۸n(�;�ջ@�~v�\gE6����Z�\��us� �����q|D[���?��Y��o��r��<ρ:��fqG����e,� �	LH�q�g��-B$����k�o�<J4:ƨ̡�nʴ5�b�!�m��ݝ,�}���e+ßBY�1�\T>)	�n�5bj�;!r�/-���t��:�^�|�����e
,g)k�{2ތ !q%�L`ECA�	y�#-�Ul��®M��̈E�V�x��
�{��u���\��jW�4ݤ4��l,>a	b�DP�j�?��v`��i�����a�^L%�;	b���Q�ӚX:��Z� �D��/�Ò�Ҷ��99��U�L���D�eK��g��܆�!��!Pk1�mX<���p7�k%jj\\0Ĳ��
�������������Y��*)Q�;�\�� ��旰�*�9�q� v}̢o��y�6l�Xv����jF������]g,��U~��V��bcq��9�iz��]�]�Tn��N�wȼ�
M�R�i�9V�s�dΦ�\/ߗ�u6��허���+��Vt� �,��%��вM�]⎻���G�[�ʹe�Iܖ`r�+�A�
?��'��[��y�<�]�B�[�ފmD�IX�-o�-����~�4���2fFO�3NOWf�5�lU/�N-*����?/�Ő��A,$H�Qp7��10���I�c�}�GQ=�Pʬ����][W�z��!��PM.������ʙXx������9ˌ���Ē�V�!妖h�nY;}��>:�â�;����d����fd���QӤgͳO��Y&GlY�-'�C��$���7�8\6�N��<WB���݀)���&&�`�l�.�D��Qf�Ƣ��OWB�d�o0*��3k�K��A:��`8Q��n��^ ǭ�� x���O%a+uZ[�*�z1.#�]{/"@�G�hĀog��n���G�OJ�������R�>F����A:_C���<o�"y��5D��5N��7M�0����c �po+��8d�����,e��X��A�yϩn�@"U��F�� ������:_���z�������<�De')����f�=�>֬�e��W�#��#i��.��Q�ߤ�Q�tϚ�l�O���T*̏L��\S�ԉ�~\�Fh;-	Iօ�c�qp��G<Ǩ����"�g��52�蝖nF��w.>�li��U�
��������9��wn�	zm\?��H������ߜ�`����O�m���|^3-��L��Fh����{��'�(6D�r��� T���s��4'��<{v��q��)�6_�e��<<_�pE�Z��7xm�z�[�m/Zq��\i�/�Z���:��ۚ���g߽�$f����F�4�1��Wթ�'��w�?��0���r�/�ǡ�b
/���ql����=�%X�ݐ����j ��|Ps�Je�#��;�Ɛ9�`2���R[�)�tm;Qo����~]�4�K�K��eA�E��F�-_���3�{ktؓ�����/W<���	g������an�De� a�n�fJ�v:����3�,�	�
��;�e�����~\p��K�a1�cyL1$& 7E��ވ��b�@/"��&Wg�D*�����t�k�}{E|]��*ŷ,r�l�\W�H��Yq��s����q#N<<<�s�~�7g[`9��tcp���B�b���氤�9ܖ/��	�TH���a+W��*��I,�a�Y���텣�KY�֣~��"���&�9��(h��#W�R�+�.��Q^c�b�H1�8��tAf2!%L���9���R���"�Y�;��+2�r�4Y<0�Wʜ�߷xP	�h����T8�����D��U���>�^��<�
>�� FTe9���*\����7	��%~���`�A��jwߨ皵gQ�tP����m��fq�,�Z��xA5X��UX���[���+�����c��>�90R�,��,�D<��u9&���ѣ!ٜ�H{Y���A�����>yzt����p��^� �c�J��� W���+�?���Y�1}���s��Ou*�����CG�y��y(\����[q����
���⦛�,��)�Ex�����I�F����x�q+Nu*L�jX	��4.��ٱ�Q��U`k_~��{��u �J�,,]��p ������ϯ|q����>�y)�k�����m�s�"ˤ}M�"�,&�;�
��,%($��y��g��,�?[NMz��3OM�8kE*�a�NI�Q'I��8�P���אE��
�&�tm��(L�
&Bg쯹�V���		6z�#��T���ޯ�")�_p����	%Ѩ��u��N�����|8��h�ݛ+��*aN�j�/wB���5Н"�r��ؤA*�O$��)�`����(` ���
*@6���}ç��y3ב�}��%is2���Y���s�����5m��9��F ���᲻�u�xj���o�EHct0���!�
�U�ڌ�
e�NL�P�r���D��=J,Q1ҳ�2P3���XA� �/�03��֗�E��!$e�9��[?w�p�0w�
 �z(Id3�� �uX_������w���3�M�nG*�d
{�Lu%ŷ�%ă�|��!��:-&�R6�/������5����LÍDF$�߬�d��k��N8���\a2��HW�m��H1��㕮_Q��j|{)��KPC�f��k6�Z'k�`�7Z�Æ-��P,�݂���#�t��$!��G˔ �_�[qo<���I�_�΀�h����;fl��Qi�&F`�PW_�ih֘�+��]����Aٽ��2ϒ#�$�F�P4�w�g\�R7�z�K[�)�8����Fv�"6Y�o&W�s-Q�l$�
��-����>o�GT��ſ���趤��L����u�N�%�S�u�~��]���N��L �V?[��:��R��s�$R����'�2�y���)�d2Э��#�'����`�N����E�*x� J����6�aར�U�s$���|8a��G
o�G3��nFS+4P�"�(Y.���Ė�C|�u��vGW*�rGS�C�ً���F�v5NY�=����t�=��
,f�R��� ���Nxv27`+�y��"��o�P�
���HǤz&�f!]'S��>ajv�$�4/��#�	,�y��[���hVP�7
>�iV�q<]�R'0e��K�$��f���w��_��FV��x��r�(Lj%����!E�/?=,�9PhY�S����;0P��������1s�=�Lv�T2�o^��h�I>p��ٲ���7��-��
Lm�h��S,�9��=��s�Iɖv�� ���jͪ��M�:s���*�B6�'y��W��o�K���p�
���$�`\i�ؗ�����A���t�>���$�v�m���������*�y?�A0��	�do	�J�>�|[���� ����}!�{���&��'�z;�$*��~֋-��hn���&��y�����>8ѻMC@� n����� ��ӁLL冞7�y���@J��3�T�ߔy��O�S��
Y���Ʈ05�J�ɀ�n�:e��qH�����:w�zp��G��w~�҄����|Gf��] {�<�U�7�45	,Fӣ��#N���2���������"g�R�ru��n��E6��m 5Q��%;h�9n,6H��fƩ�j�ۑ��v�Uճ�#�v�+�Hݓ`$�	�Ǚ7P।���vw\�Xr�-�)�=59���Ȼ9�Id�	����Z�˺�����^ as �nMIkkSrVx�x��(�y}QFo�j<ﶽA&���Ju�$S�����7����۰��A��2�/��pw_S�@=Mk^���5���2eT�}��@����:,��,�zc}��	�f�f�T/ܿ^a���r4I��|s��T��?]8~��el��S���p\hp���;�r��߰*�r6F��,e��7-�v�ڤ~�ԃ�����2�WݴZ���\_�l�/�p��-m�a��)�5�7��ؼ����F��w��j�d�U=�*��Ab���;��Z�	b�ύxÜ�~<B"�sRs_
�T�����}пhjj��3�?W^ic1��wu�^��&��S�����O���ah��ە�:��U;h�x����nFnU�e������߾�$�|��4	#���!��M.�����i���Z%�
��>O\�D޸#K�&3��t�%P���k�=M�Q�����Zѱ_܄�Bg�CC}��|��|�T ���,�F�������X��)Yn��f���`j��a���v�_غ�� lJ�� �WG_�,���� ���Y��3�TDn�t	6|ߙ�l�mْeҶ��x��G���WU/���<Q���������2@F�(��y���r�ߢ�Ҏ˳�o(4�g��!����¢%]�Ȱ�1^��1��⧟�p��)m@]�����ѵNlQ�����\=X� �8ؒ ���<R=T;��"�ˬĘHXM����5R�3��¡��@Y�i�NM޳�SZ����D��j��S��I���(��1<��C��[��v�+��"tL���
�u���F�(�m̻_z�Qc�a�^m�L.ΰԶN�~u/��,^bĂ*�4Ψ��oI�RG,�����{���Hr�dhr��u'$��p)+4�P�%��jz��9�&�S�!���XA�Ʃ��D�|��}E(#�{*e�}B�^�e)wE��ƺ9DS����)-:�/��6Q(+&��i�'"ۍ	/��
�F6
Q ̟M�a���C'T�F,�q�Igp����~�S�[��M�@x��{~�Ł�mrs��J@�g#h�CW8�O{��j��&��r��*�����ޢCó�/߀Y�{ȼd�J�qc�Oc���w�4��u*J�����n�a��!�A~�z�Qt}"Yf��;Q�PD���j��c�	��p�:z�vW��)��J�|a�=r����,���tm�E��?X�ykO��*u0ʡ�F^�<2�}bAw`�#�E�Y;5����сQ���R��g�9�}{�U4`��$��������Kv�|�:�s�$s�Χ�ۤ��Y�֣��:�ڰ+�_��gX�Q� ��T�J���I}D��᯶�9���H\�ѵƄ[�N�^+@�V3�&���ƙ���*ճܫT�f8� V�i���Ov�Z�z�t9�B�`����.LW�>'�
Ŧ|N�M��W�Ķ��>�4~ɝ�=@>��Fi'*$���c���:�w�p�%�7&j��8�(Oh���/�:18�!z�:��a<��0>�;�a�#!�WU��P�?2������r�i]���n��`��K���"������>�<5q���#x��L��f�y��A(�=���"�������P0�	��\\\�}�ƚ�p7��$�)2�r�[Ը���~a;M���B�� 9����S-��Wu�ce�s;�O��o0���kM���/l��Z��G�_Ù�K0����X̥�i��[H0��Cg�H�AN�q۷U�n\)0@ ΄�7řs��k��өw�6�9�c ���lpն�`�_�W�b�G��	��;����
�*ݑ�����Y��?'�a��Q��-��J����	?vLC+�-�_mb;a����JD|������S�a����c����ή��M{���������oiM~�H�%���"Q�Q�Y�(s��.�G�G>�)��ڶ9"�4;�>FCX�i]���2[��A�5�@�~����v�2z�2��Zc \�	+)�E�����C��of��A�b��f��)c%@��S�1+הoy̶�RrYe�������V��5����{PO&���Ʃ�E�C x�W�G-T핧��f��c�� 6z�qb��9IG��yR[�Gx&�@���<ׯ쬬�.��/)�����3�2C���������, �����	)�������\�Ww��>��Ԋ$�u��Fc���P��������u�V.�e7.��.�-����u-c�42��H��k���X�:�;� @g$R\����L�����ӭ��C����W�a��N�j^�^!Qv�V8�G���L��e�����m�x9��9��Ф�0뇆�d�P�ƈ�F��8��!V)__apѯ��)����mo�W"߸#4�(�>���]�f�����ݚZ����Y>E�
/��xӇo�� ��y���2��\�^����_�8��	���C���qK�%j�*0��P�U^f�`��n��5z��4�_}�snఞd�����乆ŢW�)�q�c���AN���33`C�X��/=.]t���.����y�����f?��LB��x�c#ݧ�z�#��������R?;�N4���Y��'��EO���%�+\wt~8���JD��~ʢRw�4F#9U��C�Vֿ=�����s����5،߆Vz0P���R1T�n1!v�6Xʈ����}فkL[�bCE �ρZ��Fvph��`����1���9(`UJ��"��W
8b�:o}���%����W6��?�H�`f�b)	&t�ϟ����P�j�&,�Y	|���+q��S*zp�kʟ��6G�Z	fA��y���+�4F	f��ψϚ+�j��|���Ls��IV,Sk��e�͎S�ڠ��s+ͣ�v��ب������Z���2�h�-- 惫dV���#�fdv�b��X��y��i�VW�J�ѯ^��c�N�p�c�2���ee4�լz(^�va�D��ED�i��Ӵt�/B�:]{V���y�eo��z8T�-�L��=G��B�@>��s3�>�љ���-�[�7�(^zv��G�x��h��,:�pg�Ý��/7�Fo�;l<�@��B��E��tw� ��Q`�7�~��l�4�4 8y:�i����2C[��V.Wٚˋǣ���o�!�� C���=6�u��#��ы������֒�)�J�]��ޘf\��"F�Q.�v�.w�2w�:�9�:[yMg5O��k�- ������L�.��B'�Ee�h �2ddc�	F�g��������z1�Ü�]��5N:����`c$��"	Wp2�k�}&�I�.&칺���6U���T�w�"�w�`y�AI:�t�[y��� H��ҽ��m�=���e�Ne�v̿����j��)�,�B6�(��&i�5���$�k̦g}�)�>�Z�%��������.��!�'�Z۹�$#?��s��do��'0p�%���;��c">EfJHs��̏�>LYJ�~�d�h�ńjIA�s���� ʬ��\�*l��3�_�K�mc�<ۤ��D��o?g�cr)m�[�!XM��\2�	d�DH�jR?'�
'i4�=`q�Ͷ�
�s�}�4��`D|��x�����}���'z�H�(���C /HĽz�q��g�¬w�~ܧh�N�k ���]��
O1�`�Ʀ����IզQ�L�c�=��X��'�{��v8�O@8��S�5�\j��Lį����!_�������'+�C[�Ow��a�'yu���Rqu���u�4D�Y� � �c
� ������1c�L��6��u���sjk	떼�K�/߃�j�Zn����|eq^�;i08bƀm��#TUT�\�����*�O�\�'I�	ͺ����c��1��r!0,���!�N���� � mD�����|�����M�g������E�������`S��v�Ě�x����E�8X�)8��łEٹU.����� c(w�RۇXYY�M�譕* �JIS����XB��k4�T'd8h��`���o~�?̸��CJ��W�_Z(E�E	���Xc���e޺yI���r�B*�?G�J���^�t�*יY�R��Z�F�V=���r�d/j-p�]��{\S���1�1�+�xNo�Mw*�"#��.H��C\\��>4T%MR��YF���R�s�Yp�:��VU�Ȓp[dVT�i�t0�56C��m�
������������y�ݻ�Vm��FmI�.ڷr~<3��d��ъ�X���B^|w/����#~��]6�U���>��qܗ��KZx2��@����c�jw���޵���{�YX̝��%b��x�i�p1?�-��^��3�Q_*��)������CJ��\.���`�w�@
������Z/�An"z���qhA�|�7Yk<�Y���q�k�|�S�ԔyUl�J��l ��M�ܲ~�ᯡ�~ĕ�����_ ��
��p @������x�Wǉ`�L ��y����(cɣ�&�+kmބݰE�8D�@ԀLƾ�o<H���pꇅ�b����$�M4����|�ڛ��3F_�I�YY�{�%�66��Η���s���opr�~�]���1�<���#�� ;"Xx������H�R�:�����F$��c�/���..z_�D���`펃(7\���VWCEL*3B88$��!~�_&� ��_�c�� ���!܄�KRYY]�g?X�����)u�p�/sZ���a�������9_E$��PL$di�K�`��é�R��U�\Cq� ���^��śƯ�5��{�F$|u�5Ҍ�NL����ӝ�:愎�%�I�DYݔ_��p�<�lŌY�������\�u;�`
ͥ��(۷��&�|�)��]f�{c9�{oBB�Z���f�:��_�٤~}�����d�F��;[a�t��
���P���r� ��	�-�9�?����=c�W:��(L͗n���մ�3�\���tG���ś`3�E,~VL �'�;gg���d<żԵv�JT4���+��u����R�>���!��#_���;;��&0���5a�����\p$���̀����<`�9�^�D��s��z�:A=��,�e�������%64�V�)S��|/�Q��x�b��`���9��5�Yi'\m�-:���U������1��］n�	l�	Zb��&�du��������dfE5��+x�Ӆ[�H�g��������(��La�u�:��=�噧����4ع�׻�����C(
6�O#Y�����bu����HD1���>=�Y���`-�������!~S����:�S�%�@��&��2E"6��Y1���5�5�ru����v$z�u7�[�rMCAa�-��2��R[Gmt튞+�z��4q��	�E$q�HM�L�O���Z���#�����T�T�~��]��;����`"x$��z��1�nُp@��ݘ��%��444���9����F��� �ɮ!����n��8���0�Uɰ�]��������h��}������U!����K6��~k�9����S�2B��e��P��£�����:U<��N������Jy�����|��-"��F*�|��"YΊ�t!���t�������*M>X�\�i�g��"�����/ɴFs����0�9��n�'+a���L	��v�t������j���񜷝���s����{6v6��oz��L0wW�^u[����S>��c��h��Y�s�����~P��Yu����9%���6�Y�l�<�g�膳.F)��i-j�Z1��eyL� ���@M*Y� �~:S丠�Q%����]
�J�R�Cӧ�0�N�l����ޡW�����E�CBB��'��g#BG�Tu_���W)��ފ���%i��
/V�^�ޅiW8οw�&'}h�"ߖ��Н�2��?n��GC�y��Jl��*�`W���v��#��ga� �C=��ټ�/H]��P����|�����^���B�W�g/�D�G}Ԩ�H^͊��L`Xg˹@��T����z)� r00��a��J|��%i�2�lx�j��E`�^{l1��}����ډ1�ܜ����YS>]�������d�z�Cp̥ d�RD;	6�a`eE��>��xF4��]=�$Ur �z���v���#��H �Y	j����^�?%��)����;����?L�K�Z�5��Ϯ��d��	����G��� i���$����WR�	:�3cp%b!}K簅��!2�g�Æ�/y�_�P��8R!?'O���F�k�����}�h�&n�������*Ҡ"���`��PJ�|y�E������ŝ="BB�'�]|%�# ���3����o���-��D�\���a��/�)�[)�كM0>hu�O_*V�ǻ�Jt�����_m!�f�Q�u���:J��NR�����\�1K��	Y���Zz�A��:��9޿`�Ͷ;� V�U5�Q�U���¤!��ώL&)�]�6��=}�X'��=m��qpWtr��4Nk=+�0�N�C+�iŬ3��AX�3��ҹ��og*DQ�h�;�=�������C C�A-�`4��*>'ܿ�p#�;�$	�M����+b��lJP#�N�������sC[�\�xv5�([K^f��%����9�Yx�F��븂_���܇Wh^T,������ld��`�3^�,%,��sٰa�����UI��pX������S���t,����H��B�H˽/���P���) ��N!���LW��0���O����i��Ɯ�>L,w�-�ʈ�p?�<EQr$nG���{ɘ�;��^mŮQ
(�X/�����+' ���M��Q�������لs�>��憎���tn��:k]�4��/���>�YEƮWI�^C�\�R��Jv$[�4�A��ݥ	�=�J��R��S���ڷ�t9$^9����c����B��G[CF3� v�T��l(.ao}4��P�G)�����J�8�u�]�����F��,�aL�<��>�{@yy-0�:%�@�P<�B������agAb�V��$*����C&�9q�YrY2W�Ϛ?^y�s����x�(@�ܑ�]���?r2��B̥3�`WOs�goD5���bs��<&�>��R�pP�2Pe�G����pG�純���.=�_kZ�^�D�@/S�Ⱦ���g�{��o��s��B���ÒBh�������֒Ȗ���@̂_:}�: -�$�A)�o�VE/E'`��Di(T��2��ϯw`KhUmm*O�������ꛜU�D�g�ӈ�t3�(<�P��r���+�D �y��b�Z �7�z2�K�+l4�@���i�+���%�+Z'��EG�f���P��o�h =��&��Y�'�ޓ��$�q��fv���2��,�	�39�ً˨�
���ٚ=�,:{a���������:�����
x9 =u�+����D�"�X"e������[ߩ���t�����n�+�p:x�wA�dy��ј��e[S�M"���8>s�Iz�&���ύq�ɳ�2�3�!�g����[+	�yN�+���xů�#�������ƻ[�(�{�^�.$��/^�_�xE��pN�f�U����+��{�z�)�M���u���S��V<�*|I
;������H���'hmO�=�r�����$�޷�ς��qO�t��J{Ӎg?x�����9����s1��0�LT}��R���~7ˍ�~��������	N��8x�2=N����<�<�p>k�)�S(-!q9#�<�׺��m�hB�c���g��*Kt�,�?��ͳ�E�Me�뤧H�M�3,�hͭ�=ؘ�,(�}�[ׄ�ܪdD���oKן��r
D��5��
5=H��Q�ӋN�[�d��N��@�����d�y�ls1v�����|��b��ڢ>�
s7�q�|�;�3Ɠ��'��i-5�$>��j����=���$t�_���l���Nͥ���b��}�1f��4/�*	��ċ��\=7_*�GXf8�bd�~9��Do����^��a�yL�����d�'�MH6�j��H;8g U&���BZ������L�O�D�zZE��{������q�G��$R�2u���Z\��Ŧ* �"!$)9ހ--8�|�z��({��b9����Ho���̍G�箳�
��)��~��fs��_[��@�t%ɷv�рQ)����	��h$WJ<+=K�C_�x�0[�j�%��<\�<�z�?�-Rͺ��]R��
�?���]��*�2�繽���m��*�)2z����+8���`=N���3�!�*�A�1l��\��8)|2ff�pвяK%u[���E�R��g���%nˡN�e6��勌��X���ݕ�8%JP�!s�|k��}���78��Y�=f�4>CI�	J��&�7э�J��P��<������4�D�Nn^5�Ҁ$�fK����"A�{�lM�/H��Ӟ�.����;;�`�*�QSX�8|��W���1�%0Yzrj�`�����"�B"�fS蟃�5�J��!r���53"}�4FV.M˅�%�`�fJ	�L1zP'�V�Sa��wVdUy.���7�0�'�Qؔo�\�bM�i'_��we���8��;two�T{�����5:�z\^=�#��=�Qs�S떔��
]#�>U~"��o��P?�]��Ib=�������m�X6���pa~�c[`#��h�&�t4_����ؐ�#)>�C/>�,r�?��/�	24Kw��� �0�d��Ƞ�
��.�&�^ҕ�PY�(�����Md�%��%y�eލ3FM#9{������ub�ux�%�!����ӹ�0��_�T������A������ظQ�Ŝfm��jv?^���f�,�^X��I,~ej��:��f]0�l�����>��-�}螝�ǒ��V�f����`e����E�Z��ʢ�k�#���b��F?q����@x��j���Wc��,]�ćüۼ�>�d���`IWt5�Ftn�y2%���[0�_�}g��h�-r��V�F�8�e){2H����*��.j�9z؂~�K�̞�����rd]�oo�"��qNξ=ݑ��I�v��~c��p���?��I)��πW��������:1�����A��5�A����������yoC��UTk�".��x�X�uf>�;#[F�k�g�v �ԕ7�?���ɰ$��t�EJ�����R�R�0B�� D	�1�Fb��ݽь�{������������u]��,r�c�-to�r`�-�+��%K��������׆nC��[ ��3JKKw�^0�e�>8	����tIC��U.iI�)0w�W�y%as����L�#O�,�,��H)6��R�sϫR*�G��;Wcuԅ��u/,�E�ȴ����Y&�;}���I��_w
w��g}u{/t�c�I�Ȁ�(���>&|`x:h�.f��Y�~w����?"l�v�qMj���.�s���R=.��p��U� �Ŝ�r*�(����;�Hoz�9�O��z_FkT�*Ro4�ғ���"�����P%��D{�l�E�A��E��" =i(o��&�ZN<`}Z���Ģ�&�����\�L遆&œ�<GE%W�e����%V�t׷o��t�/	�N�H~z�*�=�c�;��#������MлW�5{��7�����4��d�"g�O��� �3�*�t�h�+����Xzϖ����1���37�U?Z!7���.Z\H�{x�-�d����Qū��/`0���isoo�L��&��aMq�E�`uN‏����Մ��H�5ت�ŹʞF�l�h���[	�NC�(�d��P�%�~��o�$��ݽ�z���6������}��ʸ�n�\Oi�1U�5��/D���Q}X�B��2d2�E�΅��0+��.����j�������ܥ���v���q����X�����Ǜ|$qM- �'q܇�s�ta�u�'2p�Wz#7�Le��RUh���]Y)�(D��v���c[.aI��w���}f��`�7�z3p	����0�g�oD�&�0?��[J*BI
��IL�Tz5y�qC.s�颤�_�R�y��.��%��W�am�Gv��ҵ���~c��X�&G���+�{Q���c���ez8�ˎ�^[��+���1�!ɪ��h����Î� j�G�g��su�n74x���ޭ�!����l��/3fbǇ���J�tc�#-����t{ܟU�#���ٿ$e�\#���mk����rǙgEz��qD��;�OOBW�쭣7X+��dUg9��f&%�SX_�A�`���8 ;�)K���ȁ�<Wuou}O��H�z�.
5�a;o�̳�����BĦ5^S&K��nv$��h\��3�2.�NZ띒�("d��U�_/Y�����8ռ=���8�,�L�kE��&������N����t��kGG��P�W�D<o<��s�Vrk�[1^{���w~���>'�]����C�벨5�o#+��Sb�]�8�MCzl��	��i�V�k�����'+���K������9��3������WP|�&��/�땝gr]���`�[;�$;gfԸ�_���`�lR��=�FG����d�5�|9��֑ˇ� �ѹL�(�����#^k�߀�L��|$se"A0�$��=c\C~�uuą��1��ٙS�Z�/�M����rs"?�K�h���%��I��s�I�S�%��B��<j��N�AIV�E�[z�����Z�������"�;B�	dweq�|w�D��9پ�ЋYX��ż%]�۬x�y)���ꢤƷJL7w��`��{Į��`�� �,�+Y4��YY�gZ�@�T��Zaa!n��~��O����T-����|xX�7���=b�;�ڥ�h�`#�Z*�m��(��`�����N���17p�m!��Q)�q�g� R�㯏,£�ƀ�φ.�!8N0U��	���^(�m��\'�?�P���]c�h�����?\�|B����	g��ͭ�Ƨ��G��b�Ճ�y�Mw�O���y=��0"N�̫��Hk=�~]ҩ������I�;t,�cҫ�M���JiB&��H;�̕����`�a���"y�ƣg#g�k��1}�

�W�7�;ӎ��Y�͕�~0 �;��Yd��&⻯p�R��5�pq0Ѕ#^			��IW���L%��{E��z}B�.<B���cPd"C����������sq�@�9� �?T淰��b����Vt�+>K i��ȧT^���?�*+�/s�ژ��L�e)Yb9�苣�aH���ȣ��|��Pa��s��颣�J�;:v�$���t�DDg0���j;z�L�p͵��p��[���33��
@��Ą^��A�&u�������I�<ݻ����{x�g���I5�B��e��$��Ջ�<�Q���6]iR��`NH��$�J�x�����$����xjtַW��d����|���g��*ǂ4H�5E�Ip�k���ja+��&�k�G��W��`�¿�9��c�ůCD�_@��)�@���m�/ӟ�ݙA�VW�����>fD�����	<��.i퇹-ގ�P�`0X��Lq��K�g�?��R�Q��ǝK����lY�+�R{5v�aL���GHr^>7iP��L)Gb	 .�C�1��="]���:(涓o�>�I~GT���HҶb<�"J����o�:吨�����eP4$*��D��$8��R�<R@^iy�55t8��྅����$	ô7���Y���5�޼y��+nxb"�����p!΃323[��:�+�����M)�<�n�	��v\��R<���^��OK���h���j�:��Vt&��nI�b9���s�ŝ�נ�$�N�i�ެ�<��^����.�}�j:I˾^'N����z/�q0vM��y�(ztgG���$�3��n.;��2�~�vI3��	���C���ԗ%	�W����.�}o���#'�fz9�0Ш��-�ƥ��h[��;k�L���q(z2��8Z�����(u�!@ѵ�`�čj�ێ�6.?�50��b��,��uu�JD���<&��}�=��ZP���mm/z�i�����O�3N�H�`�L�݁�����	 4А���>�䥆�a�m9-P�M�+�oo�#���ԯ�)�m9b$Z��hgq���]�&)��܍g��y�O*���%s"�6�2u�a[ �a�.ۏ�e�Ɉ�������7!��s�Dh��N{��?1�[�YK��ޙ��$]dX'\�U��>�t����ר}���&tf�S�<�{�|Ձi4�L�����j9Qa�x���bp���YJ#��[�28;u��ݩ�� j����ׇ]��eŅoޜ�p͆m]c�N�'ai1I[ާRcK��� �^�����0V�L�{IZ>�q:jq]W�q�}�����N]��>�q�]
��fQ��M)ymM����.�CW��xYK�{k��^,��Y��K�}��`�����QʂH�D�����x�e	�����Prֻ�qI" S.)��>9.�Uۍe�����2�\��>p�P~\z?P4 ���t���� ��u#3�9��7�prb�G��AZ�_������H�?�?�4f��Ru�"��f��Y���￞���%$K/'���3�N3�/P�]�{�s���涤')�q��x	^��c����'}Ώ i�m�N.�,��@��A�Z�Ό35�m�[�]H�$G�r�X�0���TyE�����#1^��z$�~�ߣZT�٘�O�����G��ЯJ	0�@;�K��dK����#�&�Y�M�F��.j7n�_��P�PI�
O}{m��h<	�>�n<u����
zg�@C0}���Ks�(z����ZѪ�.&�߷�4�����3]��hd�h�k?��@�{_���ge���(�Q~��`�ԗ:s�e�C���@�
�6�_��J�i��񙮁4�������M�<�B��Q���#�p@�Їyܔ
 �Ē3Jb����H�ƞ%�5<<<��"���Pk��8J�^mRz��0"e?�J$ć��$�MEM��LD^��V�lv)�f3��V��fj�K�#p�����i}�jG��.��t�=
D�
���K���������)sF&��ϳh��^���~q�	���3����q�}�p�@[�UPPPf����\������D���o200�ʔ-3�"'�������P���p>�%M///�7TUU}��0j���e��N'|ϡ��d��¿�[�1}���@��v	����o2�=ԕ$g�ţ����gᄑ�R;���o^{�$�v%��T�DJ���6�}h8����:��7�<��؈�8�v Pꅖ�FP��钮*E>�:ύ��k��8���~��pV�Wӵ��ܱ��S�Ò��ܚ����S_�p�|[��2��/�Y����G��{���y2kx��xb����)���iӢ�������L��4�͑ۖ�7�~h�l�"�///ŝ�_d��>q�	��]����jҙ��j[Z�#X��-w�T�ۀ�&��s��"{�Do���m�Je����JU������օ|%��/r����WC^;�.�J K(��+���%����Jl��)1��������_q|zKy�Z��'nó�jl2w|w��<�,���-ǋ�b���&� �}�u��}y���c#���<��av������� �.v���ϴ�~�W~q0S>���=����k'c��߿_c�D��`Z<�Ԙ5�#q?��\snn�n`	s��n`svrx|���G�D"u��%lmm���ɳb
׃xĪ�	��u����(%��=�5�H�7U͒��˃�rv:����4Kpp(�$�����	��A�@3յ����O��@`ӕn� ��w;/�d�O�v��B�N���"�@��>~��bꍓ�#K���]K�=�w�b��}~V�ꥡ���^&4�pt�殕�nx�a��OW��:ʯ�:�$��2������i��g�d�,�>�e�b}���;���̶iY�J�^�-�
oy�!���e>�ܫ�v�9߳<��$�`k�V�?8�w��s�,���џ�'l�Q����?[���s�����{yM�	jW��d��R� �'���f�.����_��W���Z�5�\��OZ�����L�,�{�\�$y>0z��+x�ɪ���v��������`��`Y������S�5�ĚKK�(��R��{�G���3�v�:��`��7وSb��e!w�Z�V���O�{�lư[�沣���+d5��t�����/8H4v��T�E�	�+����/<rv騛D��mq����$8������ۑ􂝋�C33�11�m{��S���Z-�%j���⚛5�_�{xT���<�Y4ܫC�(P� YH6c��{�~k�.�����`#"���w�x�zw&�**�lS�o &�Iy�[�?���%{]u�r�j7j����q���-��y�񍏖�������%�&o16��Ck}@^�O;3���>��/@q�$	iA;�k����������4�ާ q��n3T¦��ۋ��$S��b�K����̪W�TGB�2�v,��oz��-�S�.=�?������H0j������O��Ĭ��s�]�㝹�o�W�n�R�؄� ǈ�zp� ���Q.����3��E����rvB��/-�����M��)©Ԇ����}r�>�'8��t%GI@�2ܒ�V��CR���ٷ��A�+�6�"�(1@|����|�����O��� q�ж���iFpI���0(�9=�?�  ���!�j�`�,R^4��``b��?Qe�^ڙ�}������]�
��(���744�y��TUW;��R%x�O������d���PܒK�^RcP?��6��h�Dk���Vdb~�q��է6��6a�h��K(dٲP�x��A?����r�OS���(]_޸8�����K��DoT����l�E*���gu>�7Rڝ!�b��X����~�䄿tO>X3=����f)��v��ɹA��˙��=�t�b�c���[�c��D��D}m��V ;�r����iX�e�g؍���##�DXn,9������D���c7ww�Ǝ��[�����C��(z����/Y{�8�=m7��f�%��wܧ�@OϚvy_,貾���릲�J�RZ�{��W�KE/�뿲����G�P<etv��$��fb�V1}(���m�R �:�L	kF9[ x5�b��psE��0��.�ʍ1�ض1Qx��!�w���܋�����q/�-1�c���9{�"��������2�&qO)f�=��S�\�<�"��m��	B�pw��XYYu�l�V���t��j$��)��cr��~Lf�s��-ҕ7����K3�Þi�!h��RE�Q��H��l7:��-���Zk
_�/�����>�Ը���A������y#���Y=�}���1��B$��鄹�L��lI �'#`�ORMԍ�
J�a�ʂ���vn��vJ�F���$��J�K��/3n��֦!��J�ɣA��$�~g��㿍@y��<��Q�7�p�5!RL��7��X�Tp�׫�|�Q�n`��ϧ�[����Ɲ��P�����v�8��W9�T(3-����m\0�OT$����r�����K.'��$?����%8�����/��Tˤ��R8�-�4�9&���o�6��A{�U�S}���T��W�0�2��N����r�O�s�_���P����^!G�?�݈�t��iQ��,�Ey�
jx0�2\i�"F!���l���/]��`��#&-��`ebaA����'��q�yW���qW,�Z�Y GFn�-��Fσ��!�`���ũ����vv|	�z55O_}n7�Y�5ITΘٹ��,�y���@�l;ۧ7�o�h��l�Ȓh9�啙k��څ�q����7�7m:#Ѻ���3��Aj�H�����uC�b!'Atx}xQ���؎�]΅��eex�MG���`�38]�iv#"u�~㾔�4_�m�X���w��[���3'V�u�O��D�3�eƿ�9$sM4kx2 4F�\�>"�pF9�x�������<j��[Y��<�Fb'��Y�4�P�#����{�cc: ��a�Y�ō@2�����w	���Qs��xx��)4��aܠP���`܍'��^-f)F�9-�YI��2 ���!�s����A��98&^�j�v�3��T,�\�vy�f�[��o@��_�y�$�(��з�]k�rB���G�g�dսl�z�an��;���x�4� Z��Ms��x*�V|�썄W�/�ˌ[�5���<�{��%j�fP�?MG�v���N�bbGǗ���^p������PiR�--�)�>LKKK��c���N����)�� j�����wB}q~I�K8\R��`���9d}=#n��ή���`hr�g;9cn`� ���pD�� ��)�J�,u������S�V�Y�VR(~gu'���W%���@K��$�y����M*�?W"�g�+�*�\"6^�Y��{.m���ʟ���fLN��b<*���o��d~M�3�p�9�����o�]��L��]p=|��K�ϴ*N�~϶�<Y���7~�$�:�~V�R?;?�j`Pbrx}!�E�&��oT��s�1���0������UT/��N�x������ַ����Xs''ʶ�6V֎�Aʐ��<EvI(555�G
4�������H���4�'aU
�RK �����ݖ���=�}�N4ų~��Na6�q#v1�v�[�zҜ�u�����S�')XR����z���r��3ukx8Ť�o(��Փ8Y#zH�ɝ��wz p.���[�1��B~+A���A�Y��3����zw㿽5H�,���������cL��fmW+�{VP�8Vvv�BQ=N5O���\��֖��߿I�ɭ��4�]]��{{�m����o��wW�_;N�7���������L��C��agg^O�<� �ITT��h[;;܏FGG�lRG�g6}e��I[t�=���S��u��|�� �A<|�4&`�nM~^>�Nà)�v�/j��04u��\:!�t����Wo�6���9����!xyZW@7���֍���b��RC�&ҹ�V4���3av�� ��s/��1~���Pwd"RT�_�u�Ay�q_���,Z�����rb�9�R����w~���n���X�	uf'��f��.��/��U�����l��{�����}a`g�g���5��͍&;;����p	?y��9a�|�㮤��p>|4!�XvNNμTMUUFv���������I�0k����W�2{Bb���5�C�w��\�C����Ip#�dP�)��������27��I���Q����i8a���%�,�Ʃ�dt���B��`|{o����ob9��>����Ǔj�I*��A�M�J��� ��Y��Z�}�j�2�_�6A�w�5/A�Z��.�`����������{��k� |��1�������T����x.�e���=3�}�n�ck������^����6�mn���S� ��/3\�q�>L[v�ل61���5��ÏO���y��B����&I4����o�����Mݐs�M�`�_�:�B��~����eT�;^�%W�}-x���0������L~�N���rCc���L���b�.Z���^��b��M?j�L}�M� }l�p����F	�c���)�|��H�Ph�8Qm���	��{��g�R���L7�O���̓;u�� ����[  �����(���v��	���\�4I����V��%t[�z�Rzy�൜��ȝp ���L}|� �V��)�231��T����K�|O��n����2X�gb�R�hV��*�1ڦЃ���TZ[k��ϖ�f���b].�Y��$���I�D���'�4%r��:OF�����GY�UR�����(7��#Z���xCf�[i2�D�^!Dhy]祊2�q�@R�0���ev��v�M��x�� "4ѧ_�wc߽�"XV��Q>�9؉Vg�Y��K�r��օȿ=�+䙠n��3���h�g z<"����-Ƈ��ڰ)�*�1b��{�6bNuk2h�ޥĜ��1�I.�.@�2[�/�17�eB���S"Ω�Z�n�;�H�آ+����W��X�U��eF����+.Z�*ff��6̍T�ۅ�$�)��cܑS{��r�i�;)��y�3�Ky����BwG�����#�i�2�Cp�i� ^�\oU�r�q(�K3E{�n�?�����"�G#s��.
�g��;�
�� S�h�mV��5�ev/v�)�eP����hR���ڃ��Q��-��gRN���G��M8��Y/qGrWGYڋ����Q���iVaֱ4����^C2ˎ��A�*��"�Ww�2��-up����,L�u0+!!x�z��B��-z�^o�*4�r�R'�9o����D�g�怯�*�}�i&��[�ۄ�\�o��������3�z	ѭ_U�M�Tl���Op��F��^Z�����LU�u�5\��_,H\,St\2�d��t8�Y!�<���3����/�������~<�?���D^�Er�d0�C�h���}��o86-_SJ(W3�0������z2�f�
�R�L��c�� KjJ�w�C�EWz^g��-K�t`k���X�N�����d G����}��"��ڦT ��?]��#�+s]��Ƥ8L��#6
��'��p{)�ݎ�j�v�]��b
3)�V�O6G���O��ud8�<���gb���fa)kM���R;�mq����-�Q8�Ӕc�>d���f��a�(�I�Zv�c�^�<`���큺�W��N�Y�2Vo#��V���뭊�3��
=	?�O����a���:ϢP��y�E�.Õ�8t�>�;��1�{�-k����-6�cAq����򞎕m�*����l��Z�Ɯf�Ŷ��!x݃G�UA(��;n�"AC�����Ût��u�"3%İ�����/�'+��j[^���&��%�]��4�����^Dl�r~Uo�r�-d��)Q�����bgI��I�1�چq�g�i/���E+nK��W_ �@ɢ�̴�z� Y�}��	��n(��=��E�%rn4L�������Փ��f�.�0�G_�8���?��O>}~1Fr9v���~��A<w#=�<�l̲�݂
�9�ŐQ�a	�tzAE�x�6G�u7L	�<��o�4N�z�9k�� �Bf+k� uիUk��z�Ս��瘸��׫eKH̦?��Y>�O��c�/BpGŠIak�w>)������8b��Χ�?��ç��� ���6	a��;4YZ���ְ�ٴ������}n��EpT��R����8(u�
���<���,��Z��`����Tʇ���9��nJ��I�C>��x.�{�*�,��8�W��X$��ίmV�#Pv��c�C��z\M�5�@f�{��\ʓdr.r?�%�U��#O�����-�6�OzRT]�&�-�i�+��O�(w���vA��z�K����[����碌��I�'�Y��Fr�-�W��[1ϳ�SM�GjȦ<��̈́s�A�"�l
4K�1���S�֒�fFj[�+l���I��R��Ty6���{e��|��3�e3��-��T%�������7<3��Ŗ&o�������>'2;���
ӱ��n#Kg*���3*�kv6��E�RyWy)G]�Rj6K�Fސxh?0���?{�JҰ%�`r|�2~�lNX��G�Z��$R�i���g��ih�0d�ȓ���IOy���0M�q�F�����eȆ\&� {ɗ�ٷ�j#��p6���0w�Mn�#�z�&!�:����,
�G�;�T��_� X��i�톇QϚ�.�@p� �8|���,�Z�v=���C�St]��. ݀]�|7F(�ܣ<�2�/ ���2���w���6�Q�܉{��Ơ��g�=ρe�<d�f�,�Na�.�\J\��4�s�|I&p2��]_EQC���1E�*�����]��EIt���I�QB���i�M�O#��eRj���}
s��>���Z;DJ���0K�(K�E�L��O���\��7�`��\��
I���8�E�=0��	G�w��|kQ����i�y���ʗ
h(��h��İ[�N�@�t	�/XH��.�����h��g�z�`��U��u�$��T�q��3BK��#g�I�`��ƩǂV�)�!q@��ئ���kN��=N�x}�sr)r��K+!���&[/�p�?��6�D�)с�,�M�f�͍U%�( �`�E���+:����`4���B���������%�zUʷW�i��in��D#)N��x�h#�uFk����x8��*ulIg���/�?���� _$�L���w�d�8����S��f&F>'�|>��ǃ;$���?��N&�
drS��~,�i�٩4j�i��o(�������	��*���/�FR����k��0��-Q\Z9+�2��q����!��3];ǵ���pD��U
�7��3�T���E�����X��|��V�W����3����{�H��-�+��tڑ�EfhB���1�D�eW�ƭ'e=gH�qI�?4���>}�}>�n�Uƛ�[�����e����]��/�M�~�����fu��׾h���Y�a���jՇ O��<f�<( X�`�zs��8N!D�,�]��>c���c�����#�b�I!�(��~�C��Q��������$<dUgV�|Wʓ�qH�%��u��GX���}�ϲP�Y�>Gꃝ8����g�4�z_L뼲H���^�x�7`V�o�*Q�!�ؘB/���8 -�nXq�Eg���c�ok/�nSu2ɸ���QC��Ee����&t�&���T%;���>8$�@gAV�=o�Gj��L��g4R*(���=���Q��k��s���u����+�<WǷ캢�袿u��:/��w�A�Ѿw&���s��nCL��޷��L�m���*��P�l�^�����(�)���%����ͬ��e9LT�4ʇpH�}x�'O�u}�e�I��S��Sy�HO��d ߬,���븡j)�}�-&�V7.(�'\�x�N�>٢{8t������k��u�>��X����La�y�RZ��TQ:�A����լ��b�l�r������Ѥҵ��I-���@���K� tAAE������'��M�@ �T��ؚt�R{�9Lk���U8�j��E6G�ף�S�Ҙsa|��C���D���P{��򩓬A�-g�-'���=u�a���}�%y�XϢC��,��s)	d&ݝ\fwYD��c�a2=��Œ#x��%�c<����g����no��ӮE����;ʻ�78���W �Y��a��}�yZ���.Y�^��7A�B�HٱST+�A�QT�1v��{��
��f_�t�Y�M�P�������.S��	yF��D�LH���޷C=��\��:��0M@�f�]ǌ�XD�p��O�@B�I7�r��<u$u��[ʾ���=�>�K���)'w<�#���6�^�cΟ��������Z��?	���F��
�&l�J�ަ��<o��i�aW�Y$�a�Iԍ�%���W[wI�;��j�D��e��V�o�o��C�7+��/��R=�~P)�����^�Za�{����KE�QY�~���l%R�P�H]X�W|�88 �4K�}{}JF�Pʭ�����p}��-6�pm�[s|�e��*j�4"��� �Ir��Ii���	9�)׈�y�M`B.��gq�z&�{����f�;uP�8�=-��"W%�}I��ӛ��s��p!�hST��5�M��Y�w�3�f9D�%�z���{<������'}Hf��|Bغ��=>��R�MN��ǡ�y2�#���+�A� k�	߄`T�)��ל�?���Gi��2\b�^��{l.�S�W{�y���ԑ�Ng��Tz+�,������ץ�Iн3/Rxޠ�q�A����=�����[֕%
|\��ꤝ&N�	7�ڦ�X2�u�o+��U�/�re5����n�i-���v=<�-��j@�Z��$�&�W�4B)�����MtȹG;�e�1���3Zyo��#��$�>�^���<v~pj�&�����_�f
�**�����6�ŭ�W��lF��^<�[z�~�xU��\�c�8=��hz������͒~�p�����&�����7�]�i��zA�l��7S�`g�U��k��,���J�Z��w�	�E[I�|M��[���S
�2WiWg�d5�Z��P���۪���[Sz*�U��l�Sޣ5�$����9P����+��,�2�}�;|���wb�AdIш��S,�m��w��N��-���\���ue<���+w�I�Q{Q�%+]W���A��Qe�w�}�@�8zv=�qjG}���w��V;j���(屖uQ)������������~�"s�ș1�6���"2�Q�{�z�$�[x�I���Gg�3�����+(�l�9i���'�s���xNɎ%�3 }��{�Ǘ�RҬ��5]W�����Yz��Ӽ�q9�=����^"JwE�-�(k�%M��#in��O��!q����q�G_��E7�CXJ��6�f��ϳ�F������vG�L�wţ��Wo�xwPՈu����G�6��p������;y�*��O׽
E!�y fl��و8cN��������N�F�����>}i�WR�JZ��@4��`��xp�C==�`u��g��E�U�Q��N�|�ƅ3ޫ�xl�+`c����x8S/�UEc��9.����� ��H�fg��L�z�!��bh.kBݡQ�/⎣{����;�L<Dm.\�X�XP�#KIZz&| ���9:c����A���&G훫�2^,+X��]f���E���ހξ�N��<Ҷ���^�
�����V_��%�<��^R� 5$�,�O&D>�m�st���Y�%�`t��W�S�P{�cC�|^�Ig���k���?8
���~z�`)���J��W��R ��^l�<����)�5c����M�;fN���/�ܧ"Dw[-�?r@/*|�It@�~G��T_��v�J�4�瞗3c|�1J4�NS�[N��W��hz���_jӱ�u?�rIe���^�6�k��o�9=��j�r�ķSK64ǉS�(P�cu�Q$Z�%ŽTmR鴢2f��K9��?�!��!A���|3Su�dō�w�7�~��oz+��~y�{H�t�<+��C�����-���q$k5�O������][ge���R�Bk|#����
�:IN�쭣��ma�{��!�~VN�Th�~%-0�ƹƴ^7/c��<o�`S+��L@��W�O�P����f1r@4jI��M��E�˸\���7F\��g�s�0%��!n�piK:!�@<�*W�:�2ڲV��Z�Dh�h�G��EhV�m险�?����%������7���CG�|
�j�A,�>���yp����S�p�����.���ڌ��Bi>��C,[����F\z�n$����
W�yD�bIhz�uӵ�ۼ��w{BA	��>׻��� s��5��c����O{��L��b�ڹ w�HRs뇹{�>��1�]'A̛��O��>��=2G]o��]naO��J�ٯ�[��&��pyd���) �.~���.����s��w�˺��e"u�7JRd���������t(;���%��zc��Vn�qd;���p}���$���#M���|)9D���|�u>ҋ���$�ն�)���<i�x�_��-/�R��Y������j�_��>�g�%�u츊a��V�uUg5�hSXDZ�"��̤�����xM@;®�d��\t=���VZ6���b��9��N��/��U/GІ���#W@~��U��z+�2Z���3c��w����`�X�@q?)Y�9%*{�hY��v��+q��>��o�3�ܢR����FW��b�!#�.���꥛�*�>G+�n�~���zf����S"�Ց��ZӛnMu�2�K{���d������0��eS�JOQ��U��e����JG�|B��d�����8�ki#�V��P��/�b�y'�HX
�vq�����������?4�W87�Aj{��'��d�w��ô�;!E'���i�)nЧ�x����m��I��%��s�NR�JV5��!�����ԙ�U3�ɹ[����[�XK��I�h}�@����%��}�6�sz�_�Lc����O;�-�(�.X;�8����9x�z9�ؚ,�2�ݿ�(��ޓ�B������4����P!oE�9�\ٰ��ii�d�������!x����Y�h5C	$b���Ч���8�&��b�p�4/�h/\҃VumNR��IU�K�\.m%�V�����1'��D��I#췜qW�ʵ�j5��/�w��'0k5��E��8zd�Oa��x� ۍg?�yI�"y�u�,���O~VV����`R�,��l��f�f�mo@���"�����l�p���_�|D�[R�4�ɨ��� |Ơ[% ��C�>GP�@=ݖ4�}�n�U_Hq���,��/�e.t�������:D�����d�$�Ąe�q�������[\����}�����k���2Jo�Df�J�ٯ���u\�=�<�����:��:n]�.88ː�8%��M�1�p��(��ϊ�Ua����=ü>����l�J4�i�7�&}�>h2}/����� ����fbd�e���ܡ��r�MHV�[>����[X'D��%��^�e���{��.U�>e��?Dy�p"�2
�B��� d�Fz,���.�TY�<ϸ;�DC���GW_J�čc�>H�Y$�$с�r
{���*P�QA�p���3���L���)����#���g�S,�y�4L�H��&7lO��HV�ũ*q����� �*&6"��$C_��R#�=nHY�}%����uB8�v� �@u������?�tB����ѺAs��f�+��^�HWj�3֏}�r�Q�E+�Dt�p8.s��q�@�c����8���x4�4qwZZ�K������)O�u~��)uL���F������� �]ze�K6���?����lw���e`�V����Њі��t�F�iq�"�_h+����:&��/��j�`ῐ����?I�P)�Պ0^�Rv�� n3X�r��o�ny�!&z��|����M�*�|��m��V�[�q#��|� 1��#���Xc���ms!��h�<>�* �:C^�)S����x7x����/t�KA!��	�(.6���i���ރF�9���ϳ�O���gL7��}�"u�'�[Ѝ�Lb�E�[�k64��?���O�j#����roX��$��o�M�㱯�w��r�H���T%p}bD�VO een������O/Y&�nr��?뎸�D��΅0�{�o�㰬_	U�Ǖ�p�ӄ�R����w�{A�ܶ��)E���jE��j�����x�ӒR�K��6��3p��*��̫�e:��\�[��3��T�bz����[�%����C|íO
�Qϐ�����b0����\2���(Y���<#>�V�8Y$��X��E����N�`�� fy�4u�x�<*��y� �!H�2�ϧ�'�W�����C�N]v)DԮg�ٙ�ѧrSN�QlfI\�"Hy�<�|��G�;����	����ra�-\�����J�S�Zw��;���-��m,xZt�`�3�ɴcJ��]��5lF=(������ʧT�R��������;�ex�
�"GO�Ai֬^�R����R���	�90�и����4���Ad#�P�Km�~ �JfXF��!)(<Uhg��P�L�ڍ�Q�kWŇ���[���N.�v3��\`.Ckn��R�������5C
>߹:0��wT����ϻ�0@�q5���~w���0O�d5��埅��ֺ%���9_���{@8g-O,1nS>sR�>��Ѕ�Ee �P���23}�:�|)��1�нO��h��Y�m}�I�l�`��
��E�Te��~�g�W����ꭣ���7P�iAT�Ni�����n$�A����CAJi�a�B������]��yך�X�����~�}�9�,_|�;vȔ]�ؽ��G�&�t�v��f�V���3^�����v,�r�xo=�-�i��һ��n?���B���B�H����@;�ү.�T�>�O��Ɇ�9�n�K�2f�$W+�*�>�	�fQ\=��R'�(�M�\I��η���v�h�<��Ag0+Zs֔hCXw�1b�?�@n�{�vv� <�y<i��ѺN�"+�!v��r�!���lk�p@��7�Q���E�k�=��ƿ��L@�H3ߌМO��FwH���^R��CN�#nn"�%wt�=����o@�-����}�k[�o5>�<���?|^^��H|��ap+�!K��2m҆�y�d�~M�Ē��+Ih�.d&��<��7���+�c�b���?G��]�
.���:��u�3�s�K3��q�dd$4]I���ϋo^=듹��}Hf�Y���?���H_ϗI"j�����`@Tc��񈅘3�M$�m�1��=���! �a@�u	f{��G�]�
R���}96���i���sQ B(���\�߈�LC��w0�7�u
 i�V��\�+�8mw:���揣�|�Ԟ��bXh!���k�=V�O�9���V��k�v�e����-�I���(Y��>6���,A���F^�����C��!���R�����'���'#�W�"+�ْ���b\�}$��d������VH���~S�b����iFş�4�h��Ӗd٣�69���.�gu��Z��D�ц��,�=�jrw��.��]cL��u4eY.�[�D4���K�+8`��wI����4ŉ�Y^�.�s���$
�K��o��}û�=?	a����50����"�
���$�!�����f��K�l�?�IВMm��F
��?���4�t��Z�-�d��.lP��{�ȖT4dg��{y�3������v�����o����R`�L&�˗R����/u$fj��-����Jɯ[�u�7�i� ����g��͡7Gh��.l��A�������߲�����Y#���S����(�����`d�-[�j�Nڑ�t'.��Vҹ������)qj�����pw1+�3���z�	΅��Byl��~���3\%qEw}��G���(���,Um-r>��BH��P&d�2����@�����8]��J����S���lw�/ڎ��H`�˳�^F���׆����������}�7j.�R�H���a����L	�vr�k��Jf��EJ�̱LŲMN�rjcz���)���. [��d���^R�K5�6ms��W�Mڴ����D��~�jmB7��(kBA��?�K`��a3�o� ��bC�L;���ܒ`�t��E����0�]D�n��}�{4� 7�#�a��ɩ%�T�!��!5�Pk�1"���)h����C�pZ^�Ʌ��p���d�OV'n��5ǋ�xOM^秵&��&���u�����X@�u�sg�>M�A`u������&�X]7�������I��r��U(�y����8-9�Qf�4<��-4�V�=��L)�%�]�xQw�H���i>�I��y�Ö%�$�W�u� ����`���
�����8y�{Q���҃U��<�̘;��sꁟG�tZѿ�����O��;6�0ި� !�;�wH�<�m4��.֬��nˣכ2~Jg`Y��@�ö
Kx���ϕ@�W:-�9U�{�1���_V�:��^КA?�j�=��$�/�1n��K��3oAZ*�QX�\�������/���J�����}��t
p*O�&�ҩ'���!0���H�ےc+8�NI�����;V�ms(F�S�r�R
h�m�zR�!H���~��ZJO���>�� �ݺ��Gǵ"��lgK�H~(������(���x�Gw��A����!�1J�sD��3j��IҬ߬�Q���U���r8O��z�^�{XR���Z���Zh��0��{�#�e����P�6o'	}�;�`/��j�yL�I	Y]�Ә�h0z�)�I�E�������x䤪�E�c�14!ݣ���n�p���(qU��9�56�t����"� A�w�������}iԢ-e�-���?2F����!^ǟ,�4U��j�l�M����^�S���V&:�V�D�����a����5H��~��v�H�LG,��>$?��,5e'�t2�N�/�m��@[����:��lk\lc�d�-��N�^����� [�<��Tv�w�g����Q��$�?�i��'J�0|����P&E������j.Y6��J�����^�J��Si�2���+� Ф�'��D|��ܹ��z���úN_ƛz���j�>A6x?��8��nxӺ���vH]� �Zv{����/�&�b���a���D-�3]#���xa��x(�3�X3`��Y����n(�$]8��;!Oֻk&G�)?yx�c=܎���?�C���wY������ag#�,��xz�M��&�QW?��%��6�J�]���w�\��(��`zu���{��y������Z�8�c����-R�Ӕ���ݔ��z����:�F�!g��!D`��&�!�(Ύ�F�#u|�; ��	�/VT	N�g��4&����Q��(ѕx�'2�3z�#ch�Q�䵼��J{
���w�mA Lg���I����J#��L�c�o���#�׾,k�Y�źq�{2�Ɂ�����z���>e��</ol�{� ��eq�t�|<��Un���T�Πz�*�ek�4��roa�mj9�\p�c]����2�W5Y�m���Dw�d���$|9g��]���/w��>�?�Ń�	]�V}�+�D���Ÿa���6���:�1Hl��'�h��@��3]c/eY�_���5��k���V$�(lA]��O/1-�����-�����b �<�����3��X5�:�:k�3ep�%5���}�ɿCn�S�;&9�ߡ��2�O��oi�6�����t����Gfp��.�[�gAa��s��������"o���_���F�<�>�gU�J�v"j����
,��d�*�R8=��k�6����g
N�^|���[�5&i�b=���z=���ƣ����X�$�	���_��Ҟ��I�~b�W�{p5�lK�ys"aruP�!?����l7&)6Ң����)"�=�7��47�~����\�����"��ގm����ZC7�ϖ�׿Nc�3�!7ߙ��e���9%U^_��ɊȄ�<ޔP�+�֟�o��S�g%I������3Z���GT(~�I}��?N�ؕ�R�?̚��栫ߨfwJ���Nt-����{�J{E1PCot&^���$��o�b1Y�n1������wx����==��X^��7O
«��9�b��6��V��}�n[z>Ps�`�Փ��l2P��J��
�J{n��@��q���ܛ�F��F�P��H���
~ .,�)�s���j1��n3�d�J1˖�*�匏m2�;b�f��V󟗺����h�������ˮ��
@�3���Y�dJ�$����t#DD��OmO�b��X�j��~�r.o#*�	giz7D\ra�������:�����������Z�F:U��ʊ���M�|�Ws���:�!w.g�Z�ۺ�
�1�)Sx���a��?h5F^ D���7�X]P��#)h������i�1^I0�$$4�dY��k�vp�>�Y�FLy��] j���W���>��=)y�q~GSL'�Gmqvt�st��"�C�����C���`	?�i6,�I��󛲪���A)C�I�>�
����eFW���i/̜=,�)�����fݬ��쾮�fP��F��b��#�^X��;=�M\������`2x�[�$���4�{#5A����������2�.I����2U=5�Ͽ����e�:� Q�ok'm=��n�_Z���pj�1 a�:U%}�Щ*�I��5�~UvD�5��|�'��G�
���OLrf���=�.����ZJP#X���b��Zyu ������{z��>	ʃ��ոG?L�G-Z�H)��i����AS�Ύ�d��C�G��dU�}�1B�|<��	N�+X#�&㉤��}K�� �\گ�_2��w��]~v��3��q��ӳ'k��yT�'[W[O�:r}7�� e�u�2y��/�.�l
@������.a}�]���Ao���n�4d�S;��*�4̝���>@pN���y`	���5r�O*����t�{y� hI��?i����$���D����n\`��=�2+��/g�^��n\aoi;~�_��Fd��^�	�G���ꄰ�p��Ə1ׁ����9r&��̺_1 Cﲢ��
&v�L(	@L.���%W�13���w>ZO���9��(DK���"7&�i@���ܿNys�fj�w ��(��g�rnd�R����8��:��������>�J ��Zh���h�Di��ӊ=T�7J�{��.�(jV�K$��!���`��������3"�.o�"~����ڤI���vlN���|�0Gz���R��:���w��00���@'�,���!g��ى�-�TI?�l�����s���O��0�:�F�����Ze���_+�q�K���WM,ڮ\�5�ׁ0:yå0���Vͳ�%��Gã��$qJ��x��]?��I� �^�_�+pt
!d�ͱH<����	�W{�3iRS�/uq���F��u���%��(SNJ
gB��-N���y+�}f}�zM�Pm�6S��n( �Ϣ���+�i*��g7�� U��d��(���/�=5� �WJ���kp5����K,I�+�׈s=?]�Ճ�z�q��qbF?���;��3)YpEk�p3B��ތMR{�:��d3�x�,?�����s�@���Z�aw�mwh=ȡ���!���V)���`Zntt-��Ώ5�fw>������o���4lm..6bBjQ��ܔa�9rt@�x�d��ۋ[wlOY3�l���5���7�
���h�Ǉ7�p�������r��?͹O]H8VO���vb����W-��L:�*�oT���0�,��W��ߘE,{5FF����<e#j���P��>�5.U-�������g����1���@�{ZMp���f\��d4٧���y>�J1/I_P�D�1z�����m�~j�H"N3�q�t>Q��ѕ��5b,Dkʄxy�ɓ���똌�#�ǡ���t��"�(�~տ:mxE�MH7��=����Qt��ѝ=͆2nD��QKɆ=�1�UKör�'��qJ���
8�Si����*t$o�s��:�~�֥N�S��4d�p�xD�A�|�}�W����W������':�E���FA	��o݅v����{~�K���z��#�(]�J��x�t��	e�P��~�B��BP��Y�9Hj7V��x6*g'���\����>�U�}��5����_���<v��סZs�ڂ�T)+L�AM�~PH��/�����u։�j��y�?��Pb�=0 �L ��G���k�������TsR�t�p��X0a'�}��4I��T�|ND<i�7��Fo��������|7�S�y��?)�$�mk��R�L��Z��)���z/S�o����8'X��G�6'�SQ2Ň�iy�ks�S��&���Ƌ�߈|�v�3��{p�x2�,Z�/s�8����b�Z�9!��\N��������:{�s���~��⹘6���2��&N�{T�Ē	��hV"�W�}���r�HV9Z�$�*��yֿ���� �Q�j��I{���z\��%H�Wx-�7�wLKV���4��8bQ�j�L�<J1rq�o��<�d�\_¥������i@�����#2���"��Jj���]a�%���ցB�Bȍ��K�E�%�/3�a��E���뎌�ж�ݻ/G�m.�yA����?� щFD%�]Z"�mda���P���"*$`<�� �;�9m|In;�1�{�5�&F�Ys�M[8��x¸���ސ�1��}z���s2ȶ)jcfQ:"�=�]~[��!��];���d������?��l��.�����*���H����a�����ݸ"����<�,��s��V�\���oO(�=¹��,)��J} q�2o�����>9�)�|BA^����cjW�xC(�æNAa_���md �_ZS�����|�j���d�|�(�=��6M��!_W�o��ۜ�a��@՞�׋�෠�bv�`�Q��_--#K���9\dt�j/U;j�Z3F���]�����o_E���A[�FQz=�&��[r.7�9�\kG
�A������:X�`��~����8�g� J qx���X�J�nb�_*0aU�m��3?_I����,s�I5ͼV�z;����^��3)�x��s�V��K� �Z��?I���.!b;���+�k�R"�w�jċ����	��I'L�)5ZT�0�F��=�Fy�����o'���������� �(SB���D�##�;T}��v~���P���̹��/�������U���&�J�^�ނ��?� �.q�Ʈ���>�)G[�ϻ����LGke���q����\�ӍSϔ#X�1�U�Xr�1�Fɱ�:`\nx_Va�b�̇��􊻲~��i�����!��(%>���o3#X��ʙ)���jז�����߄�[�wtg9U�}����.w'ؘ]����27w��(5�w�缀_7�U��O���h��a��m#���ϕ��̖qjG@��a�,����#���>���A�v�BO@L�dV�sl��º��q!��z�wI}����3l#$G,�8�{,�����o@8c3��A�?�����[�[�m�_n\�oJ�7�S�>��[�N=�!氏��iq��Z�%a�Vh�����&d�^�P�[��HF�%�f�cV��2��E�N���c��V6p/������l�a���[�/��a����������[	2�ka��k��f��;�j<s�E�}G�k�"sj�C��#��q�L7Ă���Ѱ���o��� ~QdC;L��w�f󏆍@ ���1r?r:AH�rCa�C;8�%�'�h�L�L����{*��o�@Dt�Ies���l�:�}�9�"�$h��t�NwRXZI���$�cv��ч����I�5͍��s9�B�~��m������O���I�Z&ݢ��v�U�Շm���[A	�0ha�8@���t��r�4�!6)g�L���bNyA�֝�/�s��^��ү|O�� ��L��*=�4t|��j* ���RxN*uŒ���}Q���봞*� ���v���mZ����v��ݦrM���U��f�1�����X'}��V��Eh��8Z��d��Q�Cf !���G�4��߷�`� ��R�{R=�FVv~7����|0Y��gEU���H$"ǡd�,��Cק(�74�b�듇+���>&7�IZ�MvZ��ڣ����������!�F�I'm�2Sﻡ��&�w�g�kL�I�����%X���װ �h~d�s�����H�מO�7*�a�?���YV�rw��8�����7i�s6�E �j��4���8fh)��Οz��׳s�p[����\�u�Pa;-���X	ZX�6	<�*C����H���U�	����-a+�A��H�@ta�E�n�ud ��z�=D]+�u���^<b�%��n�
\t�_ܛ�@�f����:���O�[9������-�m���su�B�TO .E:)�OIP+�G$S�����`/m-�I�r��'v͈��ڍ��� ��D]�Y�D� �Z�v��_P݀Y�cCr��g_�&�#L�8��'�>��A��oL?"gE�ť6q�N���9C����e�����ц?)���.���S�"��96f���;[vA�/�IF�����D8e-w��9���:����O~��ۋRL~g#��XO
0���i�y�RW��	�hV�ӭ
�:���{���}L����`��4�HI-ڭ�1[��օT�l�J�#�2�X�v�#��z���`B�6����D-���!Hi��ɧo�f1_r`�����U@j&M�YZ�nٳ
�'�3#
[���p��8E��bT�o��f��ƌJ����c}��O�Z�b�T��HK��E�8�N��ZA�&cu 2 ���FL6v)_GF$-�� ~D�8߿��~j���Ů>d�9����⮡8S<��3w�~=SK�	�.���Oe���X����oĽAb	H��x�J��;�N������)�ݢL��u�_d_�*x�(ĝ~�f���J�Ƚj^�N�,��Ci�o����S�#�f9UX�e<2�����`�طIe��.���x�x�<��L�iz��;�C7�g�ZN�Yo�0J�Ț�P���*Y���I�>:���ju���M����t�������|��)&�w:L1{.?����׃���J���S�_�j���il��c,�I)	��Ӝ@n'?Q�6��(�N�g��ACw�M�ly?�3wûQ�fT\�����h��T��O"y]�"��⫷�=�m�I��`�1e��m�oh�7�W��*�`���a�?��>��{Ya�6x�msSz̵V$�'�u?�;����w(�
(�hν�[s鶒D0pk>�2�j�[13�E�%1�qN�zU��Z5����U �)�Jg�K̳@�An��`�ޖ�:p~eX_Y�Q5��_�y���>kEn���&n!\�]��l���G�xU$��3*	����5��!��~U����q],B��n�釘�4�n����Jy�ދ�W��i�i�{%���J�[�,)0���Vꨇ��8�bi��8�JZj�O��&:��z��;��Y�)=΢�z8�\��f7��������\���'��I}�'�Ļ1����P`�7QL%v_�@{��{� -`N�G�0���}rϽ^4���q^9%M��]�q��ܓ�XHmPI����[�(�[�L�<���^�䮊ܓK�)�<�]-K]�߻Or%D1�')����:����;\�4���eS����`f/Zvx�B��N�����1!��B�5>���_�y��o~�\����^�.�SQ�JFT�M�#Cd�6����I�T���%N{S�A�4��C��rX+"@M���q�{'s�Dw_,n*`�?��-X���8�ͻ0�e��ۈ�ܖŉS��Kqq�8�j��l���
�à<�F�ԙ���pE�NP��I\�Waקt]��4��+��R��I4�勆.�����hN�8�~����Ĺ��I�4l���x���Z|��/��@#�W�q+�&U+t\�Y���� n�K5��jՐ�6gS��0�N�]"Џ�hգ��!vU;����i�*�0�9�c-�	��\�S�W��%�p�?�z,�8��Ҭ����W+���P<I��ȕ 4�,d�_�5 k��-Ε�i�@0��	"�OT�*[Si䜁G���j�	���%�AE-��Em���E��"O?hB��Q�.�虜v�` h�)~�ôፂ+�#
T�h�`eڭ��CV�h��C��,��,�����׬R���7d��%��?��q-�>�u����$��<)��G�;�8���H:�c/>,�+�減F�KUf�D�3�\q�_5�p,��/̕KL��zQ":�$�9�
ޖ��v��� ��tP��Pc���6	 ��>�k��C��2nj���N��T���B�=R,ع��r�*mRyk���q������¡�~�D�pt������c��f�k�Ϙr�/f�ݼ1qiH���6Y�sR��p�Y��R��i�k�[�֦��x)jS���"��A��DD�*�F(&ob\mW��ơ��e�3��"GkM�m�ŸMc���ڎA�Xn�˜�b�T����I��CF$$��9�q=O;�ݘ�I�4q�\����*�7v�Lb����)�N㵅$o ����� �NU�'��D���3Ȇf%
��Z4<��FȣL�n�R�J�mG��O�:��h]�5�y����ۦ�Ӡ�����^j?R9��ۍ@Gɦ�U[N@��Z��W��P\qY����O)~�FnJS��R��P��^�LƄBC�l��GSN��9b�(��=t��DJ$\7ǥ��y�����7���Uva0�vc��Ѻ�W�ō|���@2���Xe�h2�:ǄBbd��%ic�tZWZ��J
���ƛ�~mM)K^<��_N�jζ�_gn?y�,�$�.��dW/^�1�݉ީB��l�;���k�`٪
+���>9����O"�G�0&�5I���Gm�t4���l��"��v4��_����'T8���":�v�C��O�B�R���L6o�c��r�z�ދ��S,��'�}Wҏ'��Q�g��{I���b��t �k|�u�AS��|�_݆��_��6x�g���$����[_�kG[���i��Gw�1��\��J��K�<��*�S������R�N����z�Q��)LE���(T��~�$����G�
K�lN8����=_���|�"���ϬW���9E���2���|4Ԭ�9��ؙ~�OK�*K��F�B�D�("���T�iI#��?U�	�ԛ��w���̽]_��t`�x��^c`I�g��IK)E�L���
qA�)���]��\-�ϕ��g�Z։�\r�PM��Y7�Y�C,B���� 9	:�dϦ����9b��z��D��B2�_ўK�ܥ���D��	9�]��|h`/�}�{����T�={�9-<���%����X̽��1����|�ʅ���y޽ir�.� �цh�=�+�ɲ��^%@E���r���a�zs�wT�����͖f�;����}��c���XFt(F;p�$'`������Q���Nbt��#���Z��ױ�􎀝�\��Tk���}��'U�c	:G0W1��Z��W_ �QCU���S��E��o�#*Tæ��9�ϫv���R�ߛ�?�.����
Xǒ����-N�Q����P����\�	�r�`H�:T�v��R��'%F�iX��⽿����0}�ӗkH�#�$����4��?����͉�CF��;F];�~'��_�Zo)NG��i4]��]�ݿK��T����c� )E@��Dc�o��-�,ؕOIH" �~�;���� �7��v����h�{H?|�������6	�6�6cR$���*6D­H�ѐnŒnoBf+�2���'�&�s:Უ�%/v�}k��?�d�n�AD�O�n��̻	W:,���kY�>��k��Щʕ"�Nt�Mf���t�,�B�����0�_��k����%Xw=�o
��ί�:F�iHhTjIY�j�P�V��D�7�����}��i7��$	��A����Q}:�ɘ�Ǆ~)��dDkv�0a�?VĨ��"c
�;Q����֍��hːq��"q�:�f������m�]��(�븤�F���u��e|zx����Ӑ��;8��7�i~#Ɇ`��A��E���*Ro"���2]l�6�u��q��L�_`Σ��>��*n/,}���(Esp���w篾Ҧ�������)08�ײ������[o�b8�4^Z,�a��lP��	 ��\"�×�ĥM�hZm����,A۰mT�����4�`���E)�q�!Nr��F��0;�ٿ~}0p�8��?M�\\��X�DW��>����W�JN��*CQ��w���&k��u�`�B�L�{�����Z5���k��R��%�ũka�(�@p��A8^�%f���B�G�Q�����9��-i������>!7%j{AG�S1B�b���&��� ���|�<�]&+�7����}EF��GI�G�z�M�����V'dj�Xi�,�C�޵�˿��ތ�;߻��z	B9d:�Z!G�/��]-�\��&�xZ��F�a�H�_m2'81x��
���V�חJmp��5lI��T��\>�R}��9�c���YF���K%o��}��f)sR�u,ϒ�I9��O������ �2�8w�ܺ���~�v�`N�x�̩��^��Ǜ��|��7U��c{���O��4(-M����t����!�Q��,ȓlɞ6��qTe2Sbo65d��xC��Z�˱]K�+x��P�m�"�zF�����B+��[��k��
W�SBc��*�"�9M(M��X,#F�n *%5J� �Z :�}��7���B�UȲ�*X2%β]��b�� h���<����]3�@{˦��G��<U�&�h���p
�9c�{ڔ_����2�l6�%\EQ��3�D�J��G!����S��b��D�/ �7��3~���o��ܒ~��Ö�W�f���Ty�1� �0��B�9��R�ϔn� �sY�r�mB����gՐ ;�㍖�ΎJ����Ű���p��3��oķ��l��שk�m�J����Gof��y�l�a��מ��톖 Ŀ������g����ҷQ��&�����-�귋��+Q�gD@j`������M��<U���S+������Fj[{���G�5�o�%��ۿK�*C�$�)�Y��#V'F��A�Y ���F�%|����47)rq����j�E�\<�@V����Uh�ށ��V��Q��O��V�]��ɵ~��ܤ��3"t	��٠>׹.�qJL������|�}-����a^5��M꡵�����Ӣ��u���� /�t��'߆���Vd�zX�Aa���B����(v��=�tkuق���?�p�;���imWN�y�4(,\j�'���f�f����c�L�ɂ7�
^X�^�4�`�Avp��DF����헁���7�� ���1�>(\�ݹa�r=q���v ~3��w�&��R?K��8m\���V~c���z?��s��='
��M�_�6�;��R=��l���Oq�;�eͿߕҠ��	08��q	aR2��e�f���G�"Z�ӂ=���yfO�����%��)Ac������ʮ�������, ��9�r��I %ՠ&�O�3���Ј��'"�hco��i\�4��G�z�ZN�ݯ'(���;^�1|+�`���%����b!��Fj�SL�;���*����	�����7SNI�G�]�����bLm�IԖ<��S�S��J�ޑ����ם���mf�2�eCGA5}����g�Tk��ױ���ۻL(��*����[t[-좬�R3�:HCE8�[k��"T��2r��u{��ć��)��q�3���B]�s[����x��-���M�o�p�HH�n�o�s��ki]���՝:�x����U�谥z���%�K1o|�u}@��t��/��-�,5�A�Gѧۖ4�C����
tW�N��9�јA fo��C����:rqkNe�g���o^(1���D�cˤ�W�;�.gJ�"c�q�G�h(\n�B�Vo�.Jپ��G�]kCv�B�Ă�H�'!pGJ��d�����z\�QpK��JНᤙ��Jug�:������c�XI�UӰ	�[���e,0��!<45 �Nq���1����,����6� �"�J��V�IX��Q���)�G�ֶzz|��*:�� �aɀ�:���p/�'�I��j�$���t6U"����p"�G=cl3��܏�>\�!�n��w�o&=#ylG�n���Xw�%@(�PX�K�d_S��7ίv2ʿ���%�Hq� ���s�zɿ���9o��_�#%z\%I>W��ZF(����j�=m�K9+bM�F���,�}WhƎ(W��% x�Y��0�)���$�z����_�-��_������c�w��l-�Id���zp�n�'��k `��x�@�ߘ0��(B~i��(�j��WȔkN�4��"`ɢ!B� $i��Ì;@�����!\�|g���b��U��.O��u��+���N�Ԡ���|�u
�y���M4>M�ʆ�d�v�~�G���`h��H��p<�t?�	J�N,Bz=6��W��TqH�`~|��@�FWa�w�OS�D�	��4�4f0i�-+�f�\���RӲ])Q+�k�`�+	��>7��Z��X}�i1���˧�DbS�ʛ���_��W�(N�S�߱���%-�Q�d�ŪW�:�Zhg	������7֟��@�
�Yp~�DЕjP�׬XZ��>�z�f�zW��E`��Ί���y�����::t���p0Ư=DpH���%:��}�s���9Avh���L�a+��ٮ6n7WC� 3%��~E.�t2��\��2�� ׺G�ّA��4�����.�c�g������n!���]3N-�<W�~~&(����p��2(�0�գ~;خ5Y*�j7�ok0�6�����$�XJ� 2�y�Ibj�n�H�r�N	aO!���QV���=�Hr�t^�Qu�:�M���ӧ$�HZ��{N�]n�x	��"^xC�|��+��O�z]\}�	����?��OS`d�x:?�����d7Ͳ�,��]97E��n���C��C��:wcF9�u�hi��z؋*YK:hi1f%��ز�-��R��h*{iW"A{n��豚����xo���sRSק���5���rI��H�
�ƕ�[�zu]�W�c�\�J�/B��%�q��[�B�̗��z�X,,͛�*����ii�8����Ģ^��j�q��B.�`�1��!�۴%RT��Ê��2 ��~��KC�#��\��I<����Y���E?y��[	uX�T�.�?�3�Q����Ǆ����q9I%��5�f^�όS���M��DQ�]_T�iS��P�̷��j���WsM�5
��4�u��8󇘽�]����*iC�.��=��k.ب���Iy���:�ߠ��ݡQ�y���c���%
O5b�\�׀��/�jۍ�%�y�ߩ�a��i���S�]���Q�<@b�LC���x��I9��|�:�a~ʰ��;u�s����R`]^���PSJ�x@�������m��s�O$
+8��A��4�`��@���ʙ��ظK�s�5�Rn$�n����h~�kdУ����{��~�!3%�2!�o&��FV_ns Z������!���c����'M���� �Oh�~n,�a;_g�Z��r��Gp��oA��%#��� �~��Z����&K�;��֮쵑 S��]�y�uc��i�ӈ|�;m����j*T�z�U�2���<-H����im	1�:�g�"1Yr)Ӏ��1�-2�_)� �-E�U!O7zY.^w�/)K<����Y�]ٌ.M�F.� v��u�ѓ�[7�]�3��kɓ��u�+
c���/kq6��
����Z��;-%@�.��	Q�ֹ۠W_�!Zd�l?F;i�ƹy�U���Nb���2�_+7��}g�fp�����+p���){�f��:�Z���eX�]��|!7�(�����+�+lC�&5�y�Y0|G�X)v���v �]N��៱�(����~ƃ�Qf�A���2��)A��,��Ja��^��7i��	�)-�?9`v��'�7띾���RŊ���c�����Ԑ��}@������pj�����{x1�Y0�D1�y��):ç��d��q_Dfh�d+�^Yh�/g��A�u!2�r�M��y�V#���>�0��m����ѽ����-&�u���*��x��I�jB(Xܚ����n;dQp��sH�&����#(U��v\�4	���m���1~0��v��hw��XhN��ş��"/�_r��u/�Ē�3��b��EgM�a��dM�2,���i��X�G^B���ޝ0!Ԏ�Gz~�z�'�M�Q�D�}2�J�#FUf�80��?�xa$�~�~V).@ ��dJ����<ٶ�L�������h�{]������s��R7��쭃��pU>�ĭ�>b��1pT#^Z�EYZ9�O��y��>�{r��<s)A�q�%/M�X?B��!��3>�&�Ls���h�?�H�Cؽ���%��e_��-��!����A�7� 3�-�]Hoo���BkQ�1���S_=�(�5���g��K�2�K��ՂQ�x\��.f>��+m����wG,�/���Ŕ7_V��31�3�Ũ�*��W�5l�{�N����b����i���H%���j�e%>zز+|�f"��w��r)T��p��'2%h�74(f�_��n����J�ѕٞ<{��"��I�f���E.��fp���g������t�^J����6�a+{t|�8h_[��S.}�����7EKV�p��絯N!,Ӻ�wñ�ݕ�U�˪��3�����}��O�^��@�*L?�~�j7�����(�:���%�Y�L|vf�F.����Q�eƪ?�=+����TP�`S�\=�P���J|'��mN� ��[A.A�X�(����;��[<X������x�\���*Au��"� 4�~�16	yE�#'��:�7#�O�C��W?x����<+��f;�����S�jif�/�
��S�z	׸8ÿ�֏d�c"hɞ�ڢ��+
.��.~��NR7�z���Z�}8%bɸ����u�s��(��Ά����ej��t��/ ��ҫ��2^�(�b��^�q-�tc�P�!:O��r�@�zG��ؙ��3�~䃒zp��:&)@�[��:�LS����{����TȇEe,�Ą�w��)}������/��͟~���������}�:S��J}���$*��F�J��?d�T�]�-LKq���S�]
�P�ݡ8���-�Z�]����Z܃��~���ެ�E��9{�����<	���`� u]v5Jh���m���"Y�Y�ra��(:��d�$Ƚ	�5�7�D��M/6�x���2@���zcj���K����G)�/Ǎ�*y��#.rȲ~��S�;ώ�9��ʼ���K��@1.sD���3-(��o��`c�DА{�?d��ۯ��	"��6��-�"
;8��=Q}�^'$&�HV)���eF]d�>��������Zm�*��B��~��F�Y�9a{~��Z�������P y��8���(��MPg�D�NC>j�80�.�@cQ�^���'����4�Z,�
*�kѥ�օ���9>_�\������m*����j ��m�c��#Ǐ4w��?����N˴4q��o�\�E�Wll�jG?	7�w�"Y�w��Qَ�I�[�f\f�Ϟi�=��g�u㐈���{���f65�~�	;<�V���w��������d[&Z�ߐƔQU��4#�(-��C���4�$��j��B�Y�8���4�� s�����+o��~��W:?t�������i>�&�c�/����e?Wϴ��~=�ǝ��NbS�G����g,�~1�v���H�ڡ� �vMG`�[)����q�+��7�����Nk:��j0�5����e�G\��Z�h,ߒt��]�(F��"�y��q��V��L' �!��d�.�����3K��� 3� k�%ȣ����ꉛ<��Ȓ�⊝��>�IRO�r�<g#c�-?��P4���Y���M�9������]��l\�Ÿ,��V�x�zHL�E^�~+����B,b#䌃&�1��Y�b�E�w��y������rLxU�%k�O��*�뒄�'�MfJ��h��Or|����Y��m	^��Y����Lu8��)q3}\ߦ[V���Þ�<����a�W�5�f�sVZ�$��ݹ�CZ��w(���W1������x� ��7AT�rlT����0�q��D�P"|u�~
P�ʻ@�6�q��o��J�H��p���k�C�v���5 ���s⢤@��)\��u-���O��H�[��SϠ�Zr�!u���xH��AV	^G����!j�ԃ(!C��l����w���:��o�y s�u}���\Hһ� Qi����sѵ��y�3���)^�g�o�/�B��4�W]�����$@N[�DsW�"�
CZ��r� $)��L�<R܊���~fƴ��AK��������:��[�}��`~�4����/s��-�����40y���W������2|���Uꬌ�G�:H]$G9�Y	���W(6����59�������G����j r��a�9&�_��W�-p���-	 ���X��[����7�/QZ�����%}F�����UW���Ţ�@uڤ��v�I�^q����V-�Br����F^`l8?����(e^4��d꙼���[�h�ɡ\�����y��]"|W+����c]�8�O[J��K_�梿��߬�?�BS����mty�AR���!�d���p*���0��-I�o��uJ!�0g��n�?-
Oz 9V}zy�CD`'��ܹ�@D/�����&�u������Q�]
Z�8��#%���ܬC�VI
$n�`U�X6�M���Qx��R�ʗL�d�̻��+=�񰳤?5��K=%����IR�Q
� *W�U�>%Ѣ!��%w�)�-З2O����]00ϕ�����P8��F?�EDEX��\�>S�+���wq�^���{�pё���٠��'�S���IĞJ��ZȜ_ix������b`���Jv>:R����P�axUJ��Gc��H�4�hiE/W�������C�[�25=A9G�^BF��/~GC���c��l[����r�|`H|y�c��h���T�ʹK�:8cM�;���5)��q%�9���3b��y��y����O�2�<�6�������=�{i���f�Thm!�9ou#�Kv�E;XQ�K�aEw�nS�K��Bv7��[��6o��.{	]L���<�|Ѳ�[��)D����뷣�	��Mn���n%���*���~%gQ��},'rƶ4S.���Y�͞�[񳙗hHV+Dh�ЫΡ���x'��(��.�'��Or��a@�[�NRiI�aJ��tȂʓ����;A�<��^+�1��A�[� ���H��#D�|��%�/Cl���.�� 
�n�5���{+!�����&mA�~����
��M���a��A�o-<۹J-�
�YҖ�� ��zg%�TAp�����s'x�R<h�5l��N�3H�L���Td�R�4���˛�J��o���`��V�;E�;^�b�������ؑ���-�/"�ɱ<[��v����I�8� 1�[�&a���xS���M�ŉ��OG��TiE?!1���x���0���E�j���nR�RC35J��� �Ț�-d��;�>z���~S��c�}r�iu>a?����vo�&j��~��AÖ<W��s�_4�S��6�q���n�L��H�^V�jq�#?ycW���MƵ6T"�:,N<�^~]�e���z�J�����A[ ��لqozt�W{�_@\ ��i�^Юn��N���dwoA�����8K����&d5�Jz�oLk��F�HS�zr4����4�m��4)��Z�}r��'ѱ����_'T�^�YO�ep6��r��{��Q����|�H�NE�P��q,5]|�娂��I��8<��x�X��Q�%c=���� ���h�le=�n�S���iEp�y��p�?G�yZ���[63�vy��M;�`�z��V�d�S$Ym^�W�.����AZb�;�h�k��Ԡ��M��O���L�n	��#\ӭg�t��$�����97��Pxę"�o��v�+?� Ь*1���tYZ^���
�]�����;u�Ǯ��`aAЇ��kz��.�+2���ӄ��޻
�G�9͠��8���7��|�F���QO�0�t=��ס4��.���x����]W
�%1<��F���=��ϋ�y���5�7������+ZS=���h�X�F�<<�%��f���[w-������K�Q(���e�NK���h�u�O��G�Ztg�-R�,R�Ń���ɴ�ʜ��Jw���bsީ*цN0��/K�kN}�
��l>�Sgm�т.u�`��5�W�BM7���Փ�|n�,YZ�&��8:r�qpbIX��V��F���6��O�z;+}"��ž���	ͅ���LћV��@wu:�$�4���[��}�f�D�w��ꆖ���zF'v=7� ��e^��)A�uX�v]��Y9�ڼ�� -�t������sK竬m�aq5놪V� 6� �2b��RaI:��_o_�jW.��1�A���U�Q8�*�P��Gw���[�����w��<����)ƉWJ0k�ׯ���{IB�g� ��hgQDY�13�A����uʛ�X�e�O���W�����8�F��c(���h/g5��e����3e�H@�Tcҧ���ע�����`�JV"V��E���9���>X�Y�4S}�A�0�_h���1�)��t�[:�o�K�)�bp��&2�g|n\�VW��b���B'�KX[{�Y?t��`��zǵm���|<��Ӓ5�r/#��6Я�e�!xÕ���x�	cFef�?_�y�u��?��O�l�#�-e��� s�Џ�v��=ז�Q����T���]���H]�,�Ǯ~?���>d��
J��\�o~��hp'L
W�
��[ ��v�ť�"S��\ -�9��� �N�^ςRn��3Y��`�02�`ba���,�1��V�����к�7m%ɹ�Ի�w߱��xH�����S����"_!�)�z%�5�#���Y��l�=�3�nz�jL� D�}\X�ˌ{Y�D�+����h��8Fy��������'��լ�g4Xs�������c2�����b����z�V��@�T�?�LW�´���v/y<���G�y�=\����\�,VC���J*\���[r碫�O��"���^B��t��D"��9Ok���ɟ%V�{�*?|}�P��;���;v'���
��T��_p0GvI�z�8N]d4����뎶�J=��66j<���:.�]�]�5�8#F"M.>� *�,L�7�;FԸ��=�&$���&a�9:�;��h&��%]��B����$$����jv\��F�J'��"Ύ�����%��k�uo�)���c�g9��p׀�S�z8e�Q4l�z��>�|���pl���B�� g��i�K�Z�%�у���y�zj0����;��͇�F��u|� -�΢m�c�ݬc�Aү��5-!������Y��lӚ}��{�aE�BC��ۯ�`Z�g�ou�+�=g9v��<V�l�Eg\�ܟ������g�q��X%=P.���_����o�`�+��Ɩ�%�ሥ��F6������V[��l��nI.T��2R��U�^�eObZ���N�|�5��e���i�m��W�g�W0�*�¥x���֎o�����NY���ك/�`@>c�uc��-x|Z�F{TX��VeS�.p.���R��}0��H�L�	���n ǌ�x`�ap����%�=x]�ٕ L�x:}�+a��4m5ˢ�ÓV�=��P���
�bS�]
X�DnU�0���9�r�L����Fol<�d�[<J!��}�I��0�����g��i�{}����ϵ� �4s ��~#x�|B��v�}�����8��#�k��	�%�Fy�j�-R��T��&�KZ�t��0�����P"��kTi0ź�Ǉ8��R1�� @$�[�n8����_�C��A5g��9d�X�z�E�P�!!�{3&&p;G���.q��̑��,��q���r��R�8{b��!DȍH�i���n���#�D��L#������k)�ȵ�����#Yt�6߈�<tH4�K�ƥY��cv����vy27���\�B�&G�N$���i�/-���u��{��U�~]���U�YYl[�t��Z��|n��2u��n.�p=�6u�tR��b�ݐ��~9���B�XB���l˕
��c�4�8~;gT�S�ծ��V﷐����7�녵��F?�Bc�2=N�s��&kv6(�Nɴ���>q}����Jf�:~R�D��IX*�����/��j������f"�J8p2�\q�l��)��D��;HÌ��@��9�f�0�;`֨��o�ʁ�~"c]|��\[9��U�B��v�GǪw��?
���3�or�!L}��X"᷺�
��ȑ�ᑽ�x\��N.����fU�(;�u�M�5��ɱ"O� ��� �nHW�5d		�M�)ROC��H�k=�N]l� *���!�f�+��P>Z����RyGj۳ż��GL)'���=�{т?�ڜf�{霛y#۟�Ei�m�Y��-x���	��K���l���I;���F�;6�����������Sw[���E�X+��I_�{
״����e�:
_gAa�ʴ����^�ŅC
��;�7������� �?@�r!�]?}Ü���Z��{�sӖYJ$����R����l%���6�T�o��������#��n2���C��X�U���w�A�@�k`ےі�3�����8�:[�~��5#���j1�@�y2����f��<:���:!���K��=�L��t�$��_�;���S��\�w
��mh�h'���k@K�
y猲k{��-R�0�L#���
�RT��إ����Zx1���W���0�s��{��`h��G�V���� �����K#F����}�d"���Ƿ��+�#5�jp�FO��ij�D?#�I�TZjDmӏ雛љ7.OsR�2��36ZN;���������4|���Ѓ�T	e��`a�OX%�%{!��H���ݘ�VP 4�C4*b
pvv��!�6��HJ�k�ކ۷�a������.n��<�LMp b"���xI�4jn5|	g�)����W;û�� ��nf���Z�JZ=��� ��Ot��C	#�Y +� ˨:WA�\ �)1��ZЊL�;�[P��/"���,ū묽��Yo�F2�?��6���ـlސ��t��M�:�'���y�'Q����z�X�]׶���� ��*�����S�KN� 7�'u�{H�֪<��*sXf!mw�M��{�������[]o���ĩ�d�5o#�!��4W7,�s=~c����a��$�2[�]�~�Gn$Y�wi[o��T<�ʵ2'��h��ZW����\���.�XW��+RG�Sʾj��Y��'`����e
MS	���Q�'�i��S�Ê�X�L#�yg��(n,O�V��(X�X��F�M����JRd[�E�i�V�i<�>�8�Cz^g���ml��ث�jm�Omtp���
=�=��h��C�m�鐔�C?�]`�> $e� ��*��x��Ar�W�j*�."=�k��Gg�#U��
a��Rn������YH��M��2�m�|����E�Ғ�7�V�ңL�@�}���O� ��q+�ΣUݯ�L¦��{[�}��U�n���}�Z�s�l�t�x�yb"{.쬵�Sʋ�]��I���0
��#�����̡�q�<!F5��8����AH�֞�ۤ,ިiX��Qy�v�m6��̀:#�l��L����$��q�9��
�ء��EZQx�<c�L�g��=D����|�l�3�R��H&,�vP��U�#ױxU��݅�9�%� �f5P��p�B�\b�>�@�cɩ�X;<��w*b�����,��P�_�D�hU^4�I�y��F۱ǣ�='�%��Z�m��K������ÝЊ�C�ԟK�Y�<����艴 ��Ⱦs��D�W�d	�#����Ǿ
ܫ)Xs=�8����J��9*8��M�D��DB�*Q��f���?�˜A�eg~�4~�Rӯ� ��b��������]����o�g ���P����L�kX)�Bs��ҖM�@�o�=�h*�x��Bce�ύ�j�-ݿ���e��LU���ڢ;��������v@�cLܜ��v�S=�������f3����:m�{ߨ^ƣ�0\3�dZ��<\t�v���p/�"��P&ɘHH�s$Ij��5��9Ue(C��kM ��paVA�g�)�����w�و�+R>Mfl���NHO����v	I�n�J���+z9������~�����3�%��,�O֚��ñ���g��L�>��]5;�`җoJ����h��ҩ�Vk��D�L�P7�{ϋ�i�n���t�P��ί��?�+�������h߳'G�V)}���?���'-JW���yDR�7�ɦU��˰dbd�����#�8?�-�}.3�y3�m��d�s!�~�6!�{ϼ<*���H�r폆{���P�~��3����"����H��yՎ=}Լ� O���YB�����ϸ�&�g�(\�����6?O&�apMM�*|�1_.>(h4~��0@2r��l��h� ���ǹ��^M��`�a�ڜUv����{]H��(ה"�:w̲b��~�уmD��&�]�/���_�c��{?����:p�嫻`��~�t��SCv�"Ay��n�CA�q	c��K�ʍ�w�������B-�sI�qij��!�AZY��ݼj��܍<���XL�}4�i��G�\�F*ٚ�r��)�Еv�HW��t�(Yiw7�]����V�l^ʼ�kh����sN.
��d�u;��:����a�_M��mH���w��I)�����Yx�#��!��x!��������Oc֣{���E<��F/��^f��т��nU<iKyZF�w,�.ey_D��<�<u�0��o���b���s��Q�;���j^D�v��/�78)`�� ��h�ŏ�܍5��}4mq�TFg����1lfI52��]���J<�]O�h�X�B=�5ʪEx���<c��Y��;�6O&<����-��d��P���[c��:Yͽ�b$�z ��'�&��z�
q�����֭/	�78x�p��5*H8;4yX!���H�|X�}�cg��&g=
T7�1;�)>ݰT�\�I1��hZ Hh:ހ��a�m�l�8K#�p�x��:���C�Uy�J�� ��`���O�ΣfF�E7��NᛦW�
�~v7Q��G�LM��B��}{���U���2z�u� ?`��Og���gp��M��ώ��Eg*u0����a��(���\�u�	���	x#v�;g.:&�����a�03"���BX�����S$�F��k������-�cF�N�C��5Doy=?}������RRi��Y�Z�u� 	B��� םa@�Ml�n�LxJ�1m9�^TQp<ޢ+��jcm���`1A=��?�y�VQ��|�3��|^`��}�Td���:]&0���W�
�h C��ib�9F��X�7�¿�_(�F�=۰�[R��L;�ڼ�nC�wo�#��#��ݴ6��f���QN��M��zr��V�:��)��!�ÍD-������$�6�/�$�K<�l���:��[,���nz�~��i��Er�R�b�z��I�sFٮ�54��2���8�#�[��K	��M��%��=�b|�z�-�J�1Q��F��=U[v�8��9�zY�����t��V`/�^�W��7��ӏ&����k7i��>�T�?�I3k�^�p*���+(�$=g��9Y���c=��~�[z�U��x�d�I2��B�~��y��匓M�GFA`d.��t��:�
�s��k���v��gA�Iw��M����z��w�ܴ������'>W���5�kA�NĲ�{؈�v��c����]Gm�BE���.	�B��,Q}��ܽT>*r�BǨ!��7��u��{���'s�A<Gn�״�R��D���_L�G��y�;	eD��)��uB+1
����CcR����O�PK�7L�k��Db��� ���  H �	��ms�i+B�Sܺ�G4�Z��^Kh��D{����G�Ʋ�ݙ�ŭ3:���Y�'��Ì�`zA �>rsR,�[��������U�C�͡��i���M⟓�Ք4��X�f┻��?l�R`4�C�l12��"4�g�� �H�Yz|��k��zۮV���U�B�/�-��jPa�Ң��:�4�@��?�3C1�}�ԛlnT�L���$�|�c�ѱ��Ħ��(��
ۭVa�ed>K�O�}|���]N.n�π���^�u��m'_�@æv$�~6K�W�|؄�k���=zm�0��e�5�I)z��>]�B<u�5>g%��k.O׫��<��h\�Vn[$�\��ӣ3zO��O9�\H^n<0�����
Z�	Z�d�����o��-�py���7'q����'�O$K�RS�對�Z�0zP����Ąx͗�����5v����t���f}9F��p�t�
�)d�s���t��tqW:�g��pl����B����e|LMH��N9�1���Xd�B�l���x�Y��1G\�� �꿚��R��&���G\~}���P�\�3�@%���l�����p0�t���hZǗ�����G8b��C<�0>0�'�k��Y��'�CU�Qa��O>��|����o���M=l:^���g|M�!*��6�9��OI�%������
�?cqȐ(������o���d]o<�h��V���6=�X�1�>6^��&�{������i�*	��T�`]������������}̞���eR-�@�Y&C�{v�+�_�\#��P�Xji��m��W�V+s�6r^sW.:�kN�<��z6h�o��D�}�X�W�,�ƥfz�]�;�t)��rI�!��DI�}y�m���H(�W�{85���M�kw����=[�������w�t�dI�517��*T�!��&E��O
�Oi�d�d��������D1_ƙ���w�~"�@�y<_�w�	lw��C�yko��ޑ����o3��>��G�G=�Q�q������i�V-|�Y��Y�(ՠ�QE�8�L��f��j��zy�5������'|�)����Mv�~�C�x˒#6Z���A(�ۿ���nYs:Ʒ?�<��=�������?�::�@��Q����D�r(ֆ3b	�H�m����-i��yտ��z��ҳ�[C�f˚�3h�I� ���)��@b\P�1&�$�V��{�v���S��g/·���'��@�C/����������n&�Z�Ów.=��>g��@�R��E]��n�(#N�=' �𦇪-�3�U���ߗ��E��@w|���2���y
��|�qwF�hݨN�����OR۹L��o?J3�h���r����}�j�z��QW�}bF20������/��jI}m;�s ���z��8�����񷕞r�|�#3�0�X���@A��`I�kQL�-�����q��FPqZ~"JUGm��R���x��G��������T�=U��o�E�~�]{%�c0�C2K�7�C��=���;r����[��p��_Р�F�ƒ�o���6�-�N߼������N	�%����5���bBˤ-��.�m��_�RM��1����r[ۆ-���RJ�U�*f;�_,��7ͼr��� �i�nON��t;�Ϙ��f+��3���|�_�2����D��D��
K�� Ōg�Mѩ/�ZOs��|+����cy[H��|�����'+g�:{��!�{���w��̧�O�ZV�8%o�q�B8� �D?����l�(�K"œ���(d� �s��4zT��v�b��CPm��9.�:��ox0��u�F�+��/��׺�<�e��g�'��7�OE�	�u�>�.��\Ԝ�<[�c�ƺ�P���0N����7�2�e6{�m�����@�� ���2��t�+�\S6���E�����g�C�9�\���!ӭ��.R�Q�Ё�{�\��C���$��y��b$���>�y
C% �̩��8�g/{��+޽��m�a¯j��{�O����2D�21�p��|R�j�C������V�\
�ot�98��e �]�puC��#s�`���
*�l����r>D��͆ �f��P�\��&�k��&��]zb(�wzXp����Aْ�,���$#�*Z��B����7]t�Ǹj>Z��[�sJa���-��9Gp���uWC9�+��R¯^
5NJ@��7o�A	�n`�e����֣y�N�<��=�����菓�8#GB;��]k��G��̟�9���87R����'��Cn�����Yʀ@�X~.b����q_�}Jk���QKs!gG���2�b���D�����	���.�h�xo��s���]�u�@k�h��t�B��ѩP���WX;Q��Ȓ)I���9#yɴ�mka�us�d�ϧ���`�2-�K�'��N����T<ש����H��M�:�?&�z��|��ם�4�S��d~���d��L�I�]���V�U�9?�Cuk�Qk���b�c�%��o6W�J�o�3yC�^��Wn��^�̘�Cfq����5�}&ts�S�}��Q��9~�|��Єt�@G�ĥ��5O���,~	CUs1[9�������C�/��?���GݍV�������GK*`5]�#=_˺M���kY�\����tN���	�m
�\�x,V(����~�}#j�t�q�@C[nM"NoG���֔&q(�q�ܹ
����"�_����۸%��wfvT�[���űl�/.>���Y �u�m�����뇃�G���p7�Oe����AG�z�w�s�j�w�5?�y:� �;E]���Q����S������E�W������}]#G�ͦc%���rw�h�����a�3�S��E�[,%mݟ��,|�fE�k�h	۵;	�z���S/�W���1���s���Q)�|,5y� �E������я<[j�p˯��oOܶ���q���EDAX7N�ن�]�tuR�qi%\R8�np{W�b�Z�"�oYA�D��,J���+��;�)�F>+�&��_��s�H�w��.�N�A�}��mF���������[�UX��D���w\g�q����L���ܜ���d␳�Z��Ā	c�qϟ���o�U}������x9w���dl�h�U��z096����/+b��������4�~�)�T9:�eOSe�Pz��v:��m*@`�����(���� /*�7�I�[)��D��C"��l���j�^�����S뭐V��3���<X�xO�I�I ���k�E�֡S{���6��;�*8�?PG�>>-°��1O8�s�Ō�lG�w�XJ�.���$�I����m`US�E��M��i�@u�o]j̰>-�'����&mMu�?�VF*�գ���黺�o�s��Z����,G��2k��B�t�t����V���؝:y;���:�nd��P	%��Q������V��~;&� ���FI�����!�` �Be�[Ԕ�h�U��q��6PeF��!L���A��S7gf�H��x���?�j܈���]����_�/#wWz�t=�5]82��>n��?���L7L�ֱT�(O�]1�
/�ᦳ	��x��Y�!yV�Y/
p1�[fs����>}���s\���g���	���p/�_���*��F�AI��D��d5DְJR����:�8�Mw���/����*���e8��4��]:�1T�(�ʿ ��1�Qȡgp+F[�"��,��b� �+(�8����#ݶ�_-�e�'�j��qRE2|k��?��F���<*�j�M7�+�����z/�����NO=
1�?Y��qf�H�2��i�lRca?')�t76�\�ls���Oυ��Ѯ��4���͏)T�..z�H����W��".k����|�RSdr+ǘ���sQ�$G�B}Xtr8[#+���!Q1վc�bbk��ʫ���ӅsNg��������.�2���w�*�K�(�*�W���_��d�RF��by̵S���VX�Ge~�<|�]�xe��E2�C{�'s2�#��@���S���ja���ԑÉ��J;�?���w��g'χ�Y�ֲ���g�c�f�0Q�3�������E�V���
,q	�% ��H\;MK�:����N�|�n��D۱��;̡A[\pbU��c�]	��z����R���ޓײ�"&��K�=��g���I�4.F���$D'�</m8�k�t�i��9?��p���P6��6���%����D���f����z��֌�Q��]"Έ�ݵ/���&[���ߚF�nG5���sd�ь��z`���՜0m�E�֍?ht(Tj|�b�6�d�y������2���G݊����d��L2���?1:�#�S�k�df��m2ۛ,�#C��>�f���[i�fO�m���@�>����>���B�{�b����U}߅�E>@[.�B�Ib3��:q��'��a�fb~xjV�Z��\�T<�ΐ��a��Zl?�2O�����'�-��r��{2���>T��>|�?�¹�q6}���|. Q��P.Hn&��!�輵��f/ަ&�2P�����k��ri�ގW�D���0s+sbSr�ϔLG�O�J�8A�Q2K ~gɡr�Vۼ�	��t)�����A�j$~��#w E���{�aX;�QZ�Aڀj"��?I����Q
�Ԍ�^�hi�;��Q?M���ͪ�^iڎ�6꾝�ѤΪ4r���ic�HY�:����������x&��\�ˠ��{��z.'d��묛�f��lZ6rQ���^:�(0�O�H�	Ӻ񷽦A�$�Ug�	���KWm��`vx���z�	7x�N�}besƘ���:��M�2T�0����k�7SB���e��]$�ƶG�Ƞ2M�dR7p۟�	�G�u|TK��e�ں]�L�2�
HNSp�ۈ���+���]�U���4�tm\�DO�E�;{��@3�B<��U[7�G١�E��nTj�Tk:[g�v0Q10�jO��t΁ɼ�V82�V��O�9rk��5/PN�6�/y�N�'�*1՚�������r��Q��ɡ��e���|�֫`y���uʵ�@�T,���<�@Nt�9,��K�"{1Lrhv����h6K�.�0�Mrdq�)�p$�M2G���f�>e�Rk��/D6���Mʱ�ǟ��:�%���B���I�4�)��gQ�Ć�B'���ozKН?
P�(�_�6��Sg�L�g)=�e<�����9u�ΰSK������<������v�z2N��"�>�~���`+��5�7�ă��">J��a�#KȈ�SN�`�����1G�8���"�ƫ�Ġ�x��J���ѷ���D:�K�n7��T?먛͏r9_���b w�w5��Y��Z	�*�/�=�7._�F}��Q��]#��@��+B�d���T�������Q(�oC������K�/�柕n��Ҟ�׹����r�eS�?E�{��VH�JY�>�k��O��#��O!�ՙ�Q'���W�������tc	-�� }nz�2�9Z�����Y�Q�k��\��A���c�n8֡*������ק\��mv�r����R�X����y�_۶��Xt3��e�5i��>[B�8g���=��$���:&�s�y������>Rf�q>n׺���v4鹜�qry�=?w��n3����C���_A��?���? Q�ɪ�6a�;��j`�Ϲ���i���~3m�wb %��:�L�L���
�}��A��1�����K�C`9�O��o�@7�����=
o7��a� _P)��\���r xܿ Q"�$��>n��Sm�I��U_rf�8���{^�IJ�G繜��9�C�t-�$҅��b����W��A)5����(�!Q��?T�2��^<���#�D���=Sʻ9��m
U������K��f�S�dO̎^x>bKA&��X��O��b��`D�@G�M����{�FɌ�L? ���7,�a��6Cg�A���(Ec֍w',k�՟�,;��Wl����[tW+ �O���3љ�w���U��F���)]�]�8<��&��/���@e7�I�����Z�Zk{��v6�E���q��|�h�h����ģ��U2 �MI�:XE'�+����_�)
��aASi1�;�K+K�sy��g0�L��6ѫ�����3;h,�j>��D��<E�{�UD����q�4&�� ��l�}<���#�&q/��>ř���P
�ܩ�'Ğ�I�+6@�W[b|�FR������Z�>h��q�g�񼯇�ߝ�����b��Ɯ�^uݔ�/����g�Yb�%E^���:�R�-J��
X���Rn}��`���oC��9��ʧlE���d��K�O}��6Q�r\�9�7�+��P��포�B�ܯ���N�X��	����l�G���P(����l�J�����!�l9���H���*�\>{k�q��H��}AK��"��r+��?�Ky1������W���+XAbDc�f�#���/��J�[�bu��y�G1i�J)���
�yε7�wВL��2�����֤H���Z\Pbm�ë��-�5n��+��U)��-��6'�㐸T�Z�M�]Ƙ�_+��n|�a_��V%���6W�x!�n�*B��J��g,l��Ѡ)�k}�wCM�Cdq���Й�1�w�\|���$E��џ>9��/:8r#7P�ę�{v��f+'.���1H<��'���2g#֖�R���.��J�M�yf��>�DaASN�k�`80����L4����c���b��R�(-o�p_� ~ۙ�hL�+�g��S`������E߾�c���Im�vL(�`��{���81�N4��0"�lJp]�.!���l[��T:mE��M0`�5�\�&��mY�f��������ʡ�7�L�ۣH�:9#6��?�X"p����r������DG�cR��Vdis$��]�&*B��N�ɨ����h��K��ą�i��K��ˏ�5K��!d�e��;���=�p	Y׬UZ:�����Z �Ҧx�ꭅ8c��:#V� ��eA�y����W�k��A�;���F��'@ܦW�Jؗ�u��O&B�:��t00R?KA��6�j������!x�u���d�	�Έ�%c��d���Ʉa�~�4gjB>$J^+�x�'?H����%�C��A�ߕ��Lx���W=�_Ģ������!��\�G)"���s�T�s�����2,���PH�5$��)��4e�?����R�.W�q�j૗�~�]q�?�;B�|_��῜�}h���R�3b�̺A�|�e�+�4@�Z-��bD]b�I�������p��E�a�%�v���QM_�@�]�7���1�B����QN/�����D�.EZ��X�X^�!8\,x���|��S�<� h�G��Y+j�����|��������3�� �
�Ɗco�(f�����`K������"����l�M	�2���)��'�=�&��Jԓ#bC^*&oO �>�W��X��\��U�k?��Ά��Lř�������K]&�9R-С�&!��_���	��#�L��s��b�����lCM���%��Fd%�v,���nT+*��4{	���W#N0�>�'ę�PQzK��|gTS�ҿ�r<�*�(��4!��t� ]��@h���j����J(J=�H�R��{'t�#�����?�k�_�e��v���<�L��<��|M֡�XV�����<A��6��|�D�U���i��iH��[����-�3H����ne\��/E\�e$����?��_��}|U��v6l�VH`�5�ז1�Ӧ�ݒ�j��6�QB|�� � L.�,S#��Q�v`w!�ZI��5��U4=�&���c��J�~$k���Ti���@K���~��O�{e��sR�-��(���-�$Gzk������^�iO�;�)��DR\i]��`f���,EB��'��g�=�Uh�����V��SQ9����y�X��@,�iD: �$p�����*0E�����j�(��h0oq�2Ъ�9�����qcrw6��9�L7�&�9\���]�������(# 侽Z׫FI��9�����7?�z֏fx�֝ �0��y �����)v-np�?�yGJ�i̒�=���`���!1a7X�F�í��*���>v�'$Bs�� �����$F���-/z�THl+���ϭ�T�N�@��&�\b�-����_6G�D���=>���)�5u�_9�#>d���0A���(�/�^���j���y[�%pH��y�Y�GR� B�{�,?V��3�C��X׼�P�r c�q8ޝ������(kJ����i��VHI������hw�9�Mb�>��l�jN�Cg[�`���$��\�J�3[����D)�!�ͳ��u�����fq���1+q����8�EN$>��<�ڞ� �u��{L�_=�-G��G�F�J��iih ��7��w�
ĥ��6K���~��Y-���ě�3,1|�w��$��*qI��;�&[��j(��H�y�9S$i�S��� w7P�Ա2��&'�����}�ei�q���w�W��{Vlڃ��Hb�z��]<r�D��H����; z]�����v�>L�%:f�6�`�kޕd=1l3U�����F���9P��Ʌ��(>G�ˉ�_��+6�"*�d.S�{Z�c?��_!�,x�绶��=�hH�bJ�I��/b�����5brʯ_��R�_AN*��Ai9ֹ���x���V�ON�;������~
��l�_��=�{�׊�J/c̸�[���Q�@Y���v�(m�ܴ�RI&<|3u�2�;c?Ѝ�Ş<��~>lU����Á٣"^�Ie�9�
lC������P�#L���*�s���O�^�-}�D��H�D��S�fyhM��v#�͙��e[���h6�j�N@(�e?�?���3�;���wF1�40_\sV�joe���׉ ���}��9�{���Y�~��I^�2���/��|+�����j����ҙ��w^�1ryO���b�]Ӵb~{�|�yƺ��&�l͹����.�q����6�`<�A,����B7�$�4�1DV�H�S[�)��(}M����f_.sq���Щ�K�6���;*�]ju�'�������0&ѓ6�g��?��ҵ֍I��k���b���j��9H�0��?�}*
#�Easn&��E�'k�m��vJ�/��yu���R-L|��%JK��h�'�3L�j��:����'�P�ӧ)�p��i��ީ�%o}2�t�|>e���:h�8u�e�O��בݩ�W%~��_ݵ}gl�9�@���,V�wVP�ӌ��B���Qߟ�sA�	�3V
�}T؋L�}��H���V�5g��5i��Իb��\D�<!�ǌ�.����Q��n�k�>�_>�u+ɢ���&z�����׾4�Go�p�S��+`��j{v�FoEx�
J���a���1��ԊL���!hk���m��޼���g�e��Q����齻���%d��^�	zb��fb���_�G�s>p
�$����ck��ɬm��ú
WV��
�&G��"2O�T1~JOfW5M��ΊSc*@O��7����bؓl�12<Ŏ�0����!O%|�Q3���7ν]N~�4r�CԄ
�(���<�
��!ZI�7����E�s
�Д�ɮ/�5Cc����<DAN�:��U$���B^��	�����9ܚ�����[�1!]�A5˝�-�Ԫ���!���<)�j��2�K9�q][��ػ�+�K>s��ïK�C!G��.��db�@��#+A<֨�[������s8l�,7|��p�͛�:���񮢼��Rc;�Q g-VO���	g��ᚾl@�ȎSg�N���qP����`�-�U2(��Bxn���^�ZB���w=�I�t����8(��F�Galu�Y��\�҅ ��bP�E.��3���?.[Ⱦ��h�n��E(��6�{�U3��V���:F���U���L^���;�����>"�xD$�݈�Z�gD����n�l�p[:J����у�^���*E徕�//:s�;HK��&���ļ���yy������y�m�/��Χ�PC[Wb�猯u������H�#�g�T�y�E�Y�ce��<>W��:��5�Y�қ�"_	�����g����n����8�n�nK󕼛��*x��Ss۝ �~n!Bz�מ�6��-f[����[^�s�� eM��MǼ:��r=��@��F��s�~���j2廬�M�7��E�|&x]]'V^�����`v�>�B���I���V)�����2���I6f�l4=g��7*4a�� �>*~⺼�H�pIM6�-iFm3�����]0[��).pA�u_GAAM��P&©�T||�kH-4=�:NE��8�H
296����Z=~����^7-��u�~>����m�ys[�� ��|2���E��+O��kq㥵����b�N�V_�&�˷�r�˴S֬��ļ��ng�����WE=�\�rݼ���6�ƻX���=�|��#���K�Yd~S���{[fl��AȤi��;4��� ���Ҋ�.����Y��-�f!�e�z��������Dw��+�V�6!�>�|��xW�ڞ���B�aޜ�a=&fEҾ%�w��H�N\�
q)�s83��U���<ٵz&���:�*&C� ��I��T���wW��t8"$DY69|+M��w�辯���?7q���cZB� �ķ���F	���᧪������x�EQ]ѓMz��U)爛t�B�6N?A�ֽL�`C���w�_-��EP�3E��N�]M�H�q"D����HI{��3w�@m���jF�$�6�ZJ �B�yx��-�Vi]�O�<S�~�k��]�.�I�+���e�_v�����z��f�Q&��{(뉡p�+�s�X�����H��B����j�"5��|Zk��$�=����+=��?`4l�k��"����=3Qx4�ܘ;��Fn&]f�V���Q/D��z~գl�S]ct��ڠ~:�h�s�l�ב�Mzѵ��W<HSUiW���.��aH��O&�0U߸qRk�SM&�i-�yxńY6��˜O�5!�Y���<�(����E-��=�~��ˡ�j��a�5�����ƩU ����U�:C}vaf�Z����U�e����(�TWTjm�*���"
j]kڐ#B�Ć�V3k�^��U��wbv[�R���UҦ���b^!܄�xL)7=��<Q`!��9�9���g���&��ز���u����(l~�I��Oj:�*q�-C�x��[����d�ƅ/o�sh�
��m�C��^*���yB�b�ʑ��ؼ�`��B�\���?*��8�o�:�vU���gy�)����x"ڋ!Mc$���.��V����<�v2�mF	p�9�'�f����э,�vj
W�����5�6*�����ٻ^D�ϢۣD���&S�Pz�)vz�dy==�����2�a�5����M�:�������p���Xt6N�3G�0������c�>!�UI)z�X�~��YNs!���86�]����$UtK��3���*������6�\���+`�xU3�UQ��#=->FnU͒i�I��z�c&�҂�i=	�[�����i�ڿO�f]Ii=K1�[�D�A2b���S�]���"��
f��a�����Fs&��E�9�/�!��]&�����d�J�=����V�����>G������r1P�E�x�A��za�����(f���0*�F0^��c������l�sE�Rm�������Z�ΈL� 0�e���!�*�>�&�N�BG3#߉:���F�4�ÖP>a;�L~iɔ��u�lhk�UtWN]jdcFsT�̚e��`٧
�i��}�Hk'�'�v�)�0o��=���ꅽ� �; �5��9A%�-�3��C��!��OMY���)��՘�oÄ'M1d���j�>0�vǡ�FV����'JJ�7^�d�K��Y��Ĳ�d~Ď���t��w)����e{�l�=���w��,D�N]��V�A����Co&~2�����d�%��r%]�9�_A��RZd�yv�L�w�|Z�?��u��f�BP"(�Tm�6yS�s�,�t�!f�� �^���e.�5�ɰ�/B6MW�>#N�ڟϷ�Q��+�MNoǐ�<�p���;w)9�T��%�y�%�w�`j8c����Y�SȔI;�ku���ܪdh��'!�l�L{���F�:�<������4\��v��E,�;�݅�Cx�./�)��.�����iu�����i-6��j_�;n��g��_>re�oJX�K�27Z=�u����7m��ڊrǂ2[��:�p����id���@�D.)���o0��ZX��q� l�bTJxs5�FN�1D~;ʜ`��j_'!n��y����XH����2��qO�к;VD9��]{zr��z����T�:9����t��M�a�:����r&�I&����Q�����up�r�o̠;�x�茪r͢}���3t& �縶��Eܕ .RW�\j7#no�\a��v��E�v�yr,�˒.8��*_?ɬ��厏zsಭE�؛�ͳ���<\D�f"�<$~z��N���y��_��Ȅ��/'�
�X�ŝ��G���Ε�B7zu�����q���� ���AG=��`ŪƟN���Z}з&b�ѕ���[ZY�4� �i��Ui7��b��SB����\���O7��6�%JZܲ`�������ycD^X�90퓺%��3��@u{=4��*#3mְ>����Gh����)�Kq�f���ex��k@��r�5�2�~���"�eI���L�E	d�|#E�vee��&�����:aj�s��[q[����S^U���B�bEN�V4�v�a��\T]�3�L�߈/�jh4�H�Zv`�X�G����2�q�-��b���<����c�l��:.���L�h��N���K�x�!��2-�:P�)�$r�ʺ�)*q	�mu��XM@n0�2M��ݍK�)�\���f��y��{uP)�� +�{�d(�q�n�Y�BT�c�.�	��2<���lz�-P�}�Y�
,�P�p�j��q����	BH;�P�N_o+w��2��(�0`�d'�9�**���f�9�U�I0���@N9r��
�������7�l!6aT�9����Bp�ԟ�
@q�|�i�L�OL1Z����H��ۢ�r��3{���]��ʖƬ#��g&�DA�V+�"��{��1�	o�(_����T7����(��#���L�c����Π�O����:��hs�\+�jZS���u�����?9d/F��<�j��h���D��U�_kDܪ�v���L(E�o���5���֐�<����\�0��k_�ݔ~�o�df��|c*��&Ҵ/�t��'����+��9��:�'�eEy���.`���x;�F���0N�wI���1RW�c�W4,����	R����kgZ����D*ՙ��fɻ��c��GX:�^�͹���}BT:v���@Q��Z	��gdϣ�q�[�2����\��+�}���W�~�<j�*��N�$�@ԑo'y�!X�l�m��Ê�q�@2�5�"�����+\�E�9"�� _�#y�N�F&C��Gt}orѰ���D-�r���l��-���<����'=�P�eq���>�K\���(�S|A�7D����"$5h\�h�z>�N��?��S���ʂ��������^�$,K�Nȹ <��/Y�<˥�4r_tg��(&���I�0qd���"���i�
��g�{"�b�o���C.޷�~d��$��3����}`MG{ &�E�25����Ĉԭ��M l�����	Z�g��.ўrd�r�Ϩ�Ѻ�gg�ý#-�M����w<:�}��Q-�b\?���w�K���d��m�R��YJk(��e6��k����KxH܎^8{���3�[�i8��%×Ff꙲T"��x޺f��M���3@���$�����0h2]�G��+�#���a�v���I��Yқ���D�q��!S}'{x�ی��th�-*�ś�w����g��@�y��V��BL�e����.B ����V��"x��˜��] �+*'�a��M���*�����#���s�c�A���Ğ�~u���Y�ۼ�1��"��Q�ǂ*0�`�H6��%� ��𲎔�N�����?��ap���)��P�}��	����|-u�� ue�%��I1=j:8�~v���[�~d�T�*槣�c�EPO���X�L�n$�*4Z��o쳎o?
Q�T��|HA���ˍ�oϥ~�g�;��2q/�������\�_Ey�������P8�s�bɻ�ĝ�)�0&B(�E�z�ü+��-/?"#�E���[5a��%�}ZZ+ e"Doq�g���'Rm�U��*�����U�Gb$X	� �>�͔S;Y�`$��U祿��r <A�r2��u������#��̇9��W{���"�K`.Xfa[�U'ٜ��R��bh<��{���
R���*�* �L?>]��L:�Oy���Ot�^►1��b&(��*=G�6����2^~��s�VM������K�1�X�����|��0X��9�Ogz��@!ޜ�0IJ������M���u�}['h��ow&�_�hO�)��F�_�d��
r|k���O8ߪ����CF[�E�	�J���!��ʕ��Ǝ�/ɽ�������ukך�i���b,� ղ�pkB����?���x�tu�DЭW�PH��1'������S�R�$xxU(O|W�Ş��Db#i�����<���^,���Bo�"���HuA�2���#�i��F-YC�!���K}�.+A��P&¦�����)!'�ȡ>s�'9��ݥ�jNsO��QcC��5�eI�pO�◱�6���Q���`��	�rLaM���m�Ԁ��%��lw��Z��c)ϕ���y
L��h.7yz��Q*ɍ��S��Q��l�}�XIe��Y���ɩM ��i�e%�4�y�_���	r��LE��E��!j0���ɲ��)��S������`׆�Ǳ2ޥ������d�,��[��.�窘�J��7�߽���N#eRǢ��ɳ�8��>���	z�q0@}����j]��l�t>�)!_(VX	ݺv��V�4E[�N������3 �������$_�.��"j�����Jd6^��&�~�I���I8�H@$GT�&�bˆ�Id̲(6]����3m�[�,(,I4a������DT�k�?�\J���=��(�K%�:Y�H3�u2r}��h�׼
Q��u��m� �82"����%��L���%M�����Ċ8T��Ha}���[U�dX�>.�6+��'��tN�ʖO�ٰ�4��ƹ�NJsEa��/��~&��W�������L���zD�!�-i��1?�c7o�aR���:�SGg���pY��C+߰N��4���m����CZ'��N�I܏�_��4�i�C�"�a��Ä�$��Оqn���Yg�m��Z�̺�����'�{�V�+��f���{.M�7ʷ�G���135}^+��B�z��o��ڠ�Bo2g{�>jwb$��Q'�̐��p �7j��PX���[p��r�Aw�5e��M��W'���������b�1�n)^[F7��x ��:�����/iڰ������k�o����A-�\��Ǳ��؋�;�ͷ�pK��z/{wk�N!���V��Ҹ��u)i�x!m�������A_�F!s����?�?���_����G�/9S���ҭ'���8�������N���H1���?\��7�s?�$��_a�}T�����\b�l�255��7f��
`y^�N~��g#�m��r��|�;]mdĠ��myy�����NNN+�!��1��k+�h�����Pt��eT5���P�/���b���/��?�1m���������_�/���b���/���O���˿p��RCE[9�����PK   G��X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   G��X$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   G��X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   G��XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   G��X�C?�  -      jsons/user_defined.json�X�n�6�C@�X
�_�����@b��FA�T"t-m$m� ��g�Mi�Y��rk�͋-q��5g�}M�/ː�'�&Կ��e��,�ꦨJ��8%0Ҭ�nj���������tk�_e�wyr
�mÇ���w��+W�m]-�N�g�F��}�s�h�,)�2��g�c��)���fHgF�P��m��qu�l�An���sN���#�A����
)dp�
gU�,?���S�!��3���������eQ�y��M���a�,��A�h�XM*`�v������z���Ve�i���������P5E��b#�	<#���h��Xհ$�o���f��uyry~t�|��Ò!,�������ѯQX:��`�B�(,��I�,eWQT>DU�PES1�$��'�%���_��(œ@�`,���t�G1�3ǘ$��CZ�i�?�q�!��쟳8�RtZ��ytH(:-��":�1xF��o�#��a�q�N�i��]�iE�4�]d%Cb6���H�!��
'-16NZ:"Zr*l����RaMuD��DTGr���SPUu�1J&��8�b�LA�W:�[l"j� ���Q���#�%&����F�KND��������
ܺ��؋�7�-jhֿ�*h����Lr�(rZpę�Q�t�{�S��g,�4�˺Z��-6�a�7�u��C�=�Ͳ�l�]�zGQb�%<[�i�?V���Au��q�%������X>��x��;�؎�\�ֵ��ɽ��F���3t��*C�^��)�xc?�����yY���wg��п·���:?�|�r�ֶ���흇���GV�\�ڝ�Xf��#��)����Qe�a���,�I���L��'�%�D��rMU�e���ET�Wt�K�������<e��dF	\P����:8x���:��G�������3��D�{|Τz�����s�������~j���/����G'\�4��ϗ����U�2���Cd0�H�A׹G�S���Ad�a��/P���]�V{��~��~��۞��z�p�)��@\I(�y��&�I�[���t��(����Tj��"�F�x�\�3��<I릵u��A�J�j�0�i'ݬP���8I�I{��
<��ʇ�E`$u�;��N�G�o�샹��|wJ	�
��K�bmCr��7�g�e�?d꛷��#�$�/�������4S�6�<GD���
���x!2�%�_���o.z?r�X���������K��A5j���*X��{�0�~�S{��s,7P��Pqn82�hd-�Ya��6G�=?���ȡ���c���P �"%A;�h�Q��d
�D�|�<'2%b}~_@�vFEGDc^�/`O�?��q��d�P2��sw�*��ü=MѴ�&�m 	�rVQPPr�Y�˃B�4����s�vjCi%���$π�V3�I&�33#s�ۤ՘�KYA�nj�L�(戊�i;Rb���2"+�By:�G� ��qQ��<!�ժ��{Q_�-]ؖt���k�_>���s{X����?��X��u����i��`|u[n7���~�o"~���ϼ.����)Y����k��Y�⟺DQ����9Y�dP�O�W���6&q? >39i��='s&����=�F[�!˘ \�����GE�Q~T��qE���7PK
   G��X� �pO#  	B                  cirkitFile.jsonPK
   J��X�J �i P /             |#  images/43ea4950-057c-4494-9498-aa922855ac7b.pngPK
   J��XT��_�  K�  /             25 images/5be4124d-5fc7-4623-a6e3-e2055321e8cd.pngPK
   G��Xd��  �   /             �1 images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   G��X����H   C   /             �Q images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngPK
   G��X?S��� 2� /             �r images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   G��X��) oj /             mJ images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngPK
   G��X	��#u } /             �s images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   G��X$�8�l  �  /             G� images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   G��X$7h�!  �!  /               images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   G��XP��/�  ǽ  /             C) images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   G��X�C?�  -                �� jsons/user_defined.jsonPK      $  Y�   